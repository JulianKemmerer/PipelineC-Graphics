-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.0013417182186898273, 0.005719201933712976, 0.010096685648736121, 0.01447416936375927, 0.018851653078782414, 0.02322913679380556, 0.02760662050882871, 0.03198410422385185, 0.036361587938875006, 0.04073907165389815, 0.0451165553689213, 0.049494039083944445, 0.053871522798967585, 0.05824900651399073, 0.06262649022901388, 0.06700397394403704, 0.07138145765906019, 0.07575894137408334, 0.0801364250891065, 0.08451390880412965, 0.0888913925191528, 0.09326887623417596, 0.09764635994919911, 0.10202384366422226, 0.10640132737924542, 0.11077881109426857, 0.11515629480929174, 0.11953377852431489, 0.12391126223933802, 0.12828874595436116, 0.1326662296693843, 0.13704371338440743, 0.14142119709943057, 0.1457986808144537, 0.15017616452947685, 0.15455364824450002, 0.15893113195952316, 0.1633086156745463, 0.1676860993895694, 0.17206358310459255, 0.1764410668196157, 0.18081855053463883, 0.18519603424966197, 0.1895735179646851, 0.19395100167970825, 0.19832848539473139, 0.20270596910975452, 0.20708345282477766, 0.21146093653980083, 0.21583842025482397, 0.2202159039698471, 0.22459338768487022, 0.22897087139989336, 0.2333483551149165, 0.23772583882993964, 0.24210332254496278, 0.24648080625998595, 0.25085828997500914, 0.2552357736900323, 0.2596132574050555, 0.2639907411200786, 0.26836822483510175, 0.272745708550125, 0.27712319226514814, 0.2815006759801713, 0.2858781596951945, 0.29025564341021765, 0.29463312712524076, 0.2990106108402639, 0.30338809455528715, 0.3077655782703103, 0.3121430619853335, 0.31652054570035665, 0.3208980294153798, 0.325275513130403, 0.32965299684542615, 0.3340304805604493, 0.3384079642754725, 0.3427854479904956, 0.34716293170551876, 0.35154041542054193, 0.3559178991355651, 0.36029538285058826, 0.3646728665656115, 0.36905035028063465, 0.3734278339956578, 0.377805317710681, 0.38218280142570416, 0.3865602851407273, 0.3909377688557505, 0.39531525257077366, 0.3996927362857968, 0.40407022000081994, 0.4084477037158431, 0.41282518743086627, 0.41720267114588944, 0.4215801548609126, 0.4259576385759358, 0.430335122290959, 0.43471260600598216, 0.4390900897210053, 0.4434675734360285, 0.44784505715105166, 0.45222254086607483, 0.456600024581098, 0.46097750829612116, 0.4653549920111443, 0.46973247572616744, 0.4741099594411906, 0.4784874431562138, 0.482864926871237, 0.48724241058626017, 0.49161989430128333, 0.4959973780163065, 0.5003748617313296, 0.5047523454463527, 0.5091298291613758, 0.513507312876399, 0.5178847965914221, 0.5222622803064452, 0.5266397640214683, 0.5310172477364914, 0.5353947314515145, 0.5397722151665376, 0.5441496988815607, 0.5485271825965838, 0.552904666311607, 0.5572821500266301, 0.5616596337416532, 0.5660371174566763, 0.5704146011716994, 0.5747920848867225, 0.5791695686017456, 0.5835470523167687, 0.5879245360317918, 0.592302019746815, 0.5966795034618381, 0.6010569871768612, 0.6054344708918843, 0.6098119546069074, 0.6141894383219305, 0.6185669220369536, 0.6229444057519767, 0.6273218894669998, 0.631699373182023, 0.6360768568970461, 0.6404543406120692, 0.6448318243270923, 0.6492093080421154, 0.6535867917571385, 0.6579642754721615, 0.6623417591871846, 0.6667192429022077, 0.6710967266172309, 0.6754742103322541, 0.6798516940472772, 0.6842291777623003, 0.6886066614773234, 0.6929841451923465, 0.6973616289073696, 0.7017391126223927, 0.7061165963374159, 0.710494080052439, 0.714871563767462, 0.7192490474824851, 0.7236265311975082, 0.7280040149125313, 0.7323814986275545, 0.7367589823425776, 0.7411364660576008, 0.7455139497726239, 0.749891433487647, 0.7542689172026701, 0.7586464009176932, 0.7630238846327163, 0.7674013683477394, 0.7717788520627624, 0.7761563357777855, 0.7805338194928086, 0.7849113032078318, 0.7892887869228549, 0.7936662706378781, 0.7980437543529012, 0.8024212380679243, 0.8067987217829474, 0.8111762054979705, 0.8155536892129936, 0.8199311729280168, 0.8243086566430399, 0.8286861403580629, 0.833063624073086, 0.8374411077881091, 0.8418185915031322, 0.8461960752181553, 0.8505735589331784, 0.8549510426482017, 0.8593285263632248, 0.8637060100782479, 0.868083493793271, 0.8724609775082941, 0.8768384612233172, 0.8812159449383403, 0.8855934286533633, 0.8899709123683864, 0.8943483960834095, 0.8987258797984327, 0.9031033635134558, 0.9074808472284789, 0.9118583309435021, 0.9162358146585252, 0.9206132983735483, 0.9249907820885714, 0.9293682658035946, 0.9337457495186177, 0.9381232332336408, 0.9425007169486638, 0.9468782006636869, 0.95125568437871, 0.9556331680937331, 0.9600106518087562, 0.9643881355237793, 0.9687656192388024, 0.9731431029538257, 0.9775205866688488, 0.9818980703838719, 0.986275554098895, 0.9906530378139181, 0.9950305215289412, 0.9994080052439642]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 42
entity render_pixel_368CLK_a505fdde is
port(
 clk : in std_logic;
 global_to_module : in render_pixel_global_to_module_t;
 i : in unsigned(15 downto 0);
 j : in unsigned(15 downto 0);
 return_output : out pixel_t);
end render_pixel_368CLK_a505fdde;
architecture arch of render_pixel_368CLK_a505fdde is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 368;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
signal COMB_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
-- Stage 1
signal REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal REG_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
signal REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
signal COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal COMB_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
signal COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
-- Stage 2
signal REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal REG_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
signal REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
signal COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal COMB_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
signal COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
-- Stage 3
signal REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
signal COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
-- Stage 4
signal REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
signal COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
-- Stage 5
signal REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
signal COMB_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal COMB_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
-- Stage 6
-- Stage 7
signal REG_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 8
signal REG_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 9
signal REG_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 10
signal REG_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 11
signal REG_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 12
signal REG_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 13
signal REG_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 14
signal REG_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 15
signal REG_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 16
signal REG_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 17
signal REG_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 18
signal REG_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 19
signal REG_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 20
signal REG_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 21
signal REG_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 22
signal REG_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 23
signal REG_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 24
signal REG_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 25
signal REG_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 26
signal REG_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 27
signal REG_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 28
signal REG_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 29
signal REG_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 30
signal REG_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 31
signal REG_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 32
signal REG_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 33
signal REG_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 34
signal REG_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 35
signal REG_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 36
signal REG_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 37
signal REG_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 38
signal REG_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 39
signal REG_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 40
signal REG_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 41
signal REG_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 42
signal REG_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 43
signal REG_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 44
signal REG_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 45
signal REG_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 46
signal REG_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 47
signal REG_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 48
signal REG_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 49
signal REG_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 50
signal REG_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 51
signal REG_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 52
signal REG_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 53
signal REG_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 54
signal REG_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 55
signal REG_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 56
signal REG_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 57
signal REG_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 58
signal REG_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 59
signal REG_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 60
signal REG_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 61
signal REG_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 62
signal REG_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 63
signal REG_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 64
signal REG_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 65
signal REG_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 66
signal REG_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 67
signal REG_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 68
signal REG_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 69
signal REG_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 70
signal REG_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 71
signal REG_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 72
signal REG_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 73
signal REG_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 74
signal REG_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 75
signal REG_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 76
signal REG_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 77
signal REG_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 78
signal REG_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 79
signal REG_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 80
signal REG_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 81
signal REG_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 82
signal REG_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 83
signal REG_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 84
signal REG_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 85
signal REG_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 86
signal REG_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 87
signal REG_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 88
signal REG_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 89
signal REG_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 90
signal REG_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 91
signal REG_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 92
signal REG_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 93
signal REG_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 94
signal REG_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 95
signal REG_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 96
signal REG_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 97
signal REG_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 98
signal REG_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 99
signal REG_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 100
signal REG_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 101
signal REG_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 102
signal REG_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 103
signal REG_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 104
signal REG_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 105
signal REG_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 106
signal REG_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 107
signal REG_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 108
signal REG_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 109
signal REG_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 110
signal REG_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 111
signal REG_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 112
signal REG_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 113
signal REG_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 114
signal REG_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 115
signal REG_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 116
signal REG_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 117
signal REG_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 118
signal REG_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 119
signal REG_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 120
signal REG_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 121
signal REG_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 122
signal REG_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 123
signal REG_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 124
signal REG_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 125
signal REG_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 126
signal REG_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 127
signal REG_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 128
signal REG_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 129
signal REG_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 130
signal REG_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 131
signal REG_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 132
signal REG_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 133
signal REG_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 134
signal REG_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 135
signal REG_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 136
signal REG_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 137
signal REG_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 138
signal REG_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 139
signal REG_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 140
signal REG_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 141
signal REG_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 142
signal REG_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 143
signal REG_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 144
signal REG_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 145
signal REG_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 146
signal REG_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 147
signal REG_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 148
signal REG_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 149
signal REG_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 150
signal REG_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 151
signal REG_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 152
signal REG_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 153
signal REG_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 154
signal REG_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 155
signal REG_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 156
signal REG_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 157
signal REG_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 158
signal REG_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 159
signal REG_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 160
signal REG_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 161
signal REG_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 162
signal REG_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 163
signal REG_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 164
signal REG_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 165
signal REG_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 166
signal REG_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 167
signal REG_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 168
signal REG_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 169
signal REG_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 170
signal REG_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 171
signal REG_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 172
signal REG_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 173
signal REG_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 174
signal REG_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 175
signal REG_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 176
signal REG_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 177
signal REG_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 178
signal REG_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 179
signal REG_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 180
signal REG_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 181
signal REG_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 182
signal REG_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 183
signal REG_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 184
signal REG_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 185
signal REG_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 186
signal REG_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 187
signal REG_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 188
signal REG_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 189
signal REG_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 190
signal REG_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 191
signal REG_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 192
signal REG_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 193
signal REG_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 194
signal REG_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 195
signal REG_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 196
signal REG_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 197
signal REG_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 198
signal REG_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 199
signal REG_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 200
signal REG_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 201
signal REG_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 202
signal REG_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 203
signal REG_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 204
signal REG_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 205
signal REG_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 206
signal REG_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 207
signal REG_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 208
signal REG_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 209
signal REG_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 210
signal REG_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 211
signal REG_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 212
signal REG_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 213
signal REG_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 214
signal REG_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 215
signal REG_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 216
signal REG_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 217
signal REG_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 218
signal REG_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 219
signal REG_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 220
signal REG_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 221
signal REG_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 222
signal REG_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 223
signal REG_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 224
signal REG_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 225
signal REG_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 226
signal REG_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 227
signal REG_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 228
signal REG_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 229
signal REG_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 230
signal REG_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 231
signal REG_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 232
signal REG_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 233
signal REG_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 234
signal REG_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 235
signal REG_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 236
signal REG_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 237
signal REG_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 238
signal REG_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 239
signal REG_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 240
signal REG_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 241
signal REG_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 242
signal REG_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 243
signal REG_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 244
signal REG_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 245
signal REG_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 246
signal REG_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 247
signal REG_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 248
signal REG_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 249
signal REG_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 250
signal REG_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 251
signal REG_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 252
signal REG_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 253
signal REG_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 254
signal REG_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 255
signal REG_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 256
signal REG_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 257
signal REG_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 258
signal REG_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 259
signal REG_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 260
signal REG_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 261
signal REG_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 262
signal REG_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 263
signal REG_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 264
signal REG_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 265
signal REG_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 266
signal REG_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 267
signal REG_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 268
signal REG_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 269
signal REG_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 270
signal REG_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 271
signal REG_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 272
signal REG_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 273
signal REG_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 274
signal REG_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 275
signal REG_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 276
signal REG_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 277
signal REG_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 278
signal REG_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 279
signal REG_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 280
signal REG_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 281
signal REG_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 282
signal REG_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 283
signal REG_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 284
signal REG_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 285
signal REG_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 286
signal REG_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 287
signal REG_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 288
signal REG_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 289
signal REG_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 290
signal REG_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 291
signal REG_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 292
signal REG_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 293
signal REG_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 294
signal REG_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 295
signal REG_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 296
signal REG_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 297
signal REG_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 298
signal REG_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 299
signal REG_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 300
signal REG_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 301
signal REG_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 302
signal REG_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 303
signal REG_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 304
signal REG_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 305
signal REG_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 306
signal REG_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 307
signal REG_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 308
signal REG_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 309
signal REG_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 310
signal REG_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 311
signal REG_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 312
signal REG_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 313
signal REG_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 314
signal REG_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 315
signal REG_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 316
signal REG_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 317
signal REG_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 318
signal REG_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 319
signal REG_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 320
signal REG_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 321
signal REG_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 322
signal REG_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 323
signal REG_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 324
signal REG_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 325
signal REG_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 326
signal REG_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 327
signal REG_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 328
signal REG_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 329
signal REG_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 330
signal REG_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 331
signal REG_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 332
signal REG_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 333
signal REG_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 334
signal REG_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 335
signal REG_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 336
signal REG_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 337
signal REG_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 338
signal REG_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 339
signal REG_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 340
signal REG_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 341
signal REG_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 342
signal REG_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 343
signal REG_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 344
signal REG_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 345
signal REG_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 346
signal REG_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 347
signal REG_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 348
signal REG_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 349
signal REG_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 350
signal REG_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 351
signal REG_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 352
signal REG_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 353
signal REG_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 354
signal REG_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 355
signal REG_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 356
signal REG_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 357
signal REG_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 358
signal REG_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 359
signal REG_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 360
signal REG_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 361
signal REG_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 362
signal REG_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 363
signal REG_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 364
signal REG_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 365
signal REG_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
-- Stage 366
signal REG_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal REG_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse : unsigned(7 downto 0);
signal REG_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse : unsigned(7 downto 0);
signal REG_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse : unsigned(7 downto 0);
signal COMB_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal COMB_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse : unsigned(7 downto 0);
signal COMB_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse : unsigned(7 downto 0);
signal COMB_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse : unsigned(7 downto 0);
-- Stage 367
-- Each function instance gets signals
-- CONST_SL_1[tr_pipelinec_gen_c_l530_c16_86ea]
signal CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_x : signed(15 downto 0);
signal CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output : signed(15 downto 0);

-- BIN_OP_MINUS[tr_pipelinec_gen_c_l531_c8_94ad]
signal BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_left : signed(15 downto 0);
signal BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_right : signed(12 downto 0);
signal BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output : signed(16 downto 0);

-- CONST_SL_1[tr_pipelinec_gen_c_l532_c16_046d]
signal CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_x : signed(15 downto 0);
signal CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output : signed(15 downto 0);

-- BIN_OP_MINUS[tr_pipelinec_gen_c_l533_c9_4b79]
signal BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_left : signed(12 downto 0);
signal BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_right : signed(15 downto 0);
signal BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output : signed(16 downto 0);

-- fixed_make_from_short[tr_pipelinec_gen_c_l538_c33_b52e]
signal fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_a : signed(15 downto 0);
signal fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output : fixed;

-- fixed_shr[tr_pipelinec_gen_c_l538_c23_82ce]
signal fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_a : fixed;
signal fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_shift : signed(5 downto 0);
signal fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output : fixed;

-- fixed_make_from_double[tr_pipelinec_gen_c_l538_c70_46cc]
signal fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_a : std_logic_vector(22 downto 0);
signal fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output : fixed;

-- fixed_mul[tr_pipelinec_gen_c_l538_c13_ffb3]
signal fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_left : fixed;
signal fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_right : fixed;
signal fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output : fixed;

-- fixed_make_from_short[tr_pipelinec_gen_c_l539_c33_31d5]
signal fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_a : signed(15 downto 0);
signal fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output : fixed;

-- fixed_shr[tr_pipelinec_gen_c_l539_c23_7550]
signal fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_a : fixed;
signal fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_shift : signed(5 downto 0);
signal fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output : fixed;

-- fixed_make_from_double[tr_pipelinec_gen_c_l539_c70_69e8]
signal fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_a : std_logic_vector(22 downto 0);
signal fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output : fixed;

-- fixed_mul[tr_pipelinec_gen_c_l539_c13_9a90]
signal fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_left : fixed;
signal fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_right : fixed;
signal fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output : fixed;

-- BIN_OP_INFERRED_MULT[tr_pipelinec_gen_c_l542_c24_cc3d]
signal BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_left : unsigned(22 downto 0);
signal BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_right : unsigned(15 downto 0);
signal BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output : unsigned(38 downto 0);

-- CONST_SR_11[tr_pipelinec_gen_c_l542_c24_cb53]
signal CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_x : unsigned(38 downto 0);
signal CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output : unsigned(38 downto 0);

-- BIN_OP_GTE[tr_pipelinec_gen_c_l544_c12_1c23]
signal BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_left : unsigned(15 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_right : unsigned(3 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output : unsigned(0 downto 0);

-- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c12_5895]
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_left : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_right : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[tr_pipelinec_gen_c_l544_c33_633d]
signal BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_left : unsigned(3 downto 0);
signal BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_right : unsigned(15 downto 0);
signal BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output : unsigned(16 downto 0);

-- BIN_OP_LT[tr_pipelinec_gen_c_l544_c29_d00f]
signal BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
signal BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_right : unsigned(16 downto 0);
signal BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output : unsigned(0 downto 0);

-- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c29_766f]
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_left : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_right : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[tr_pipelinec_gen_c_l544_c12_48d6]
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_right : unsigned(0 downto 0);
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output : unsigned(0 downto 0);

-- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c12_ae4d]
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_left : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_right : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output : unsigned(0 downto 0);

-- BIN_OP_GT[tr_pipelinec_gen_c_l544_c61_d9c5]
signal BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_left : unsigned(15 downto 0);
signal BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_right : unsigned(3 downto 0);
signal BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output : unsigned(0 downto 0);

-- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c61_beb7]
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_left : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_right : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[tr_pipelinec_gen_c_l544_c12_925a]
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_left : unsigned(0 downto 0);
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output : unsigned(0 downto 0);

-- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c12_6cb4]
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_left : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_right : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output : unsigned(0 downto 0);

-- BIN_OP_LT[tr_pipelinec_gen_c_l544_c82_eedf]
signal BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_left : unsigned(15 downto 0);
signal BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_right : unsigned(5 downto 0);
signal BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output : unsigned(0 downto 0);

-- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c82_478a]
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_left : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_right : unsigned(0 downto 0);
signal BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[tr_pipelinec_gen_c_l544_c12_d8f8]
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_left : unsigned(0 downto 0);
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
signal BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output : unsigned(0 downto 0);

-- pix_b_MUX[tr_pipelinec_gen_c_l544_c3_e881]
signal pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue : unsigned(7 downto 0);
signal pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse : unsigned(7 downto 0);
signal pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output : unsigned(7 downto 0);

-- pix_g_MUX[tr_pipelinec_gen_c_l544_c3_e881]
signal pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue : unsigned(7 downto 0);
signal pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse : unsigned(7 downto 0);
signal pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output : unsigned(7 downto 0);

-- pix_r_MUX[tr_pipelinec_gen_c_l544_c3_e881]
signal pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
signal pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue : unsigned(7 downto 0);
signal pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse : unsigned(7 downto 0);
signal pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output : unsigned(7 downto 0);

-- render_pixel_internal[tr_pipelinec_gen_c_l550_c16_85da]
signal render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_x : fixed;
signal render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_y : fixed;
signal render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output : fixed3;

-- CONST_SR_2[tr_pipelinec_gen_c_l551_c20_29b3]
signal CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_x : signed(21 downto 0);
signal CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output : signed(21 downto 0);

-- CONST_SR_2[tr_pipelinec_gen_c_l552_c20_c1b4]
signal CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_x : signed(21 downto 0);
signal CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output : signed(21 downto 0);

-- CONST_SR_2[tr_pipelinec_gen_c_l553_c20_6ab8]
signal CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_x : signed(21 downto 0);
signal CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output : signed(21 downto 0);

-- BIN_OP_GTE[tr_pipelinec_gen_c_l554_c14_8e81]
signal BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_left : unsigned(15 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_right : unsigned(8 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output : unsigned(0 downto 0);

-- MUX[tr_pipelinec_gen_c_l554_c14_f66a]
signal MUX_tr_pipelinec_gen_c_l554_c14_f66a_cond : unsigned(0 downto 0);
signal MUX_tr_pipelinec_gen_c_l554_c14_f66a_iftrue : unsigned(7 downto 0);
signal MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse : unsigned(7 downto 0);
signal MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output : unsigned(7 downto 0);

-- BIN_OP_GTE[tr_pipelinec_gen_c_l555_c14_77f4]
signal BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_left : unsigned(15 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_right : unsigned(8 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output : unsigned(0 downto 0);

-- MUX[tr_pipelinec_gen_c_l555_c14_6d28]
signal MUX_tr_pipelinec_gen_c_l555_c14_6d28_cond : unsigned(0 downto 0);
signal MUX_tr_pipelinec_gen_c_l555_c14_6d28_iftrue : unsigned(7 downto 0);
signal MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse : unsigned(7 downto 0);
signal MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output : unsigned(7 downto 0);

-- BIN_OP_GTE[tr_pipelinec_gen_c_l556_c14_374a]
signal BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_left : unsigned(15 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_right : unsigned(8 downto 0);
signal BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output : unsigned(0 downto 0);

-- MUX[tr_pipelinec_gen_c_l556_c14_02b9]
signal MUX_tr_pipelinec_gen_c_l556_c14_02b9_cond : unsigned(0 downto 0);
signal MUX_tr_pipelinec_gen_c_l556_c14_02b9_iftrue : unsigned(7 downto 0);
signal MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse : unsigned(7 downto 0);
signal MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output : unsigned(7 downto 0);

function CONST_REF_RD_pixel_t_pixel_t_787c( ref_toks_0 : pixel_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned) return pixel_t is
 
  variable base : pixel_t; 
  variable return_output : pixel_t;
begin
      base := ref_toks_0;
      base.b := ref_toks_1;
      base.g := ref_toks_2;
      base.r := ref_toks_3;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea
CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea : entity work.CONST_SL_1_int16_t_0CLK_de264c78 port map (
CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_x,
CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output);

-- BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad
BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad : entity work.BIN_OP_MINUS_int16_t_int13_t_1CLK_c9fe58b1 port map (
clk,
BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_left,
BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_right,
BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output);

-- CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d
CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d : entity work.CONST_SL_1_int16_t_0CLK_de264c78 port map (
CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_x,
CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output);

-- BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79
BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79 : entity work.BIN_OP_MINUS_int13_t_int16_t_1CLK_c9fe58b1 port map (
clk,
BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_left,
BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_right,
BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output);

-- fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e
fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e : entity work.fixed_make_from_short_0CLK_23f04728 port map (
fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_a,
fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output);

-- fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce
fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce : entity work.fixed_shr_0CLK_6a3d4cae port map (
fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_a,
fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_shift,
fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output);

-- fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc
fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc : entity work.fixed_make_from_double_0CLK_38477f9e port map (
fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_a,
fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output);

-- fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3
fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3 : entity work.fixed_mul_5CLK_70b28c19 port map (
clk,
fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_left,
fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_right,
fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output);

-- fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5
fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5 : entity work.fixed_make_from_short_0CLK_23f04728 port map (
fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_a,
fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output);

-- fixed_shr_tr_pipelinec_gen_c_l539_c23_7550
fixed_shr_tr_pipelinec_gen_c_l539_c23_7550 : entity work.fixed_shr_0CLK_6a3d4cae port map (
fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_a,
fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_shift,
fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output);

-- fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8
fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8 : entity work.fixed_make_from_double_0CLK_38477f9e port map (
fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_a,
fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output);

-- fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90
fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90 : entity work.fixed_mul_5CLK_70b28c19 port map (
clk,
fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_left,
fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_right,
fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output);

-- BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d
BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d : entity work.BIN_OP_INFERRED_MULT_uint23_t_uint16_t_2CLK_d9e4e3ca port map (
clk,
BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_left,
BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_right,
BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output);

-- CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53
CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53 : entity work.CONST_SR_11_uint39_t_0CLK_de264c78 port map (
CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_x,
CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output);

-- BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23
BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23 : entity work.BIN_OP_GTE_uint16_t_uint4_t_1CLK_52497a46 port map (
clk,
BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_left,
BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_right,
BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output);

-- BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895 : entity work.BIN_OP_NEQ_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_left,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_right,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output);

-- BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d
BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d : entity work.BIN_OP_PLUS_uint4_t_uint16_t_1CLK_ab623c35 port map (
clk,
BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_left,
BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_right,
BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output);

-- BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f
BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f : entity work.BIN_OP_LT_uint16_t_uint17_t_1CLK_8ed726ba port map (
clk,
BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left,
BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_right,
BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output);

-- BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f : entity work.BIN_OP_NEQ_uint1_t_uint1_t_1CLK_541f6485 port map (
clk,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_left,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_right,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output);

-- BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_right,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output);

-- BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d : entity work.BIN_OP_NEQ_uint1_t_uint1_t_1CLK_ceb57ac8 port map (
clk,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_left,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_right,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output);

-- BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5
BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5 : entity work.BIN_OP_GT_uint16_t_uint4_t_1CLK_52497a46 port map (
clk,
BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_left,
BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_right,
BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output);

-- BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7 : entity work.BIN_OP_NEQ_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_left,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_right,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output);

-- BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_left,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output);

-- BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4 : entity work.BIN_OP_NEQ_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_left,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_right,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output);

-- BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf
BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf : entity work.BIN_OP_LT_uint16_t_uint6_t_1CLK_52497a46 port map (
clk,
BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_left,
BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_right,
BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output);

-- BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a : entity work.BIN_OP_NEQ_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_left,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_right,
BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output);

-- BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8 : entity work.BIN_OP_AND_uint1_t_uint1_t_1CLK_0dcc764a port map (
clk,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_left,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right,
BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output);

-- pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881
pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881 : entity work.MUX_uint1_t_uint8_t_uint8_t_1CLK_a9a2737d port map (
clk,
pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue,
pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse,
pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output);

-- pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881
pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881 : entity work.MUX_uint1_t_uint8_t_uint8_t_1CLK_a9a2737d port map (
clk,
pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue,
pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse,
pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output);

-- pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881
pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881 : entity work.MUX_uint1_t_uint8_t_uint8_t_1CLK_a9a2737d port map (
clk,
pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue,
pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse,
pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output);

-- render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da
render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da : entity work.render_pixel_internal_360CLK_987815b4 port map (
clk,
global_to_module.render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da,
render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_x,
render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_y,
render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output);

-- CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3
CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3 : entity work.CONST_SR_2_int22_t_0CLK_de264c78 port map (
CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_x,
CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output);

-- CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4
CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4 : entity work.CONST_SR_2_int22_t_0CLK_de264c78 port map (
CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_x,
CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output);

-- CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8
CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8 : entity work.CONST_SR_2_int22_t_0CLK_de264c78 port map (
CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_x,
CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output);

-- BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81
BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81 : entity work.BIN_OP_GTE_uint16_t_uint9_t_1CLK_c580f7b9 port map (
clk,
BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_left,
BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_right,
BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output);

-- MUX_tr_pipelinec_gen_c_l554_c14_f66a
MUX_tr_pipelinec_gen_c_l554_c14_f66a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_tr_pipelinec_gen_c_l554_c14_f66a_cond,
MUX_tr_pipelinec_gen_c_l554_c14_f66a_iftrue,
MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse,
MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output);

-- BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4
BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4 : entity work.BIN_OP_GTE_uint16_t_uint9_t_1CLK_c580f7b9 port map (
clk,
BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_left,
BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_right,
BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output);

-- MUX_tr_pipelinec_gen_c_l555_c14_6d28
MUX_tr_pipelinec_gen_c_l555_c14_6d28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_tr_pipelinec_gen_c_l555_c14_6d28_cond,
MUX_tr_pipelinec_gen_c_l555_c14_6d28_iftrue,
MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse,
MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output);

-- BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a
BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a : entity work.BIN_OP_GTE_uint16_t_uint9_t_1CLK_c580f7b9 port map (
clk,
BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_left,
BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_right,
BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output);

-- MUX_tr_pipelinec_gen_c_l556_c14_02b9
MUX_tr_pipelinec_gen_c_l556_c14_02b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_tr_pipelinec_gen_c_l556_c14_02b9_cond,
MUX_tr_pipelinec_gen_c_l556_c14_02b9_iftrue,
MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse,
MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 i,
 j,
 -- Registers
 -- Stage 0
 REG_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left,
 -- Stage 1
 REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left,
 REG_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left,
 REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right,
 REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right,
 -- Stage 2
 REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left,
 REG_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left,
 REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right,
 REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right,
 -- Stage 3
 REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left,
 REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right,
 REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right,
 -- Stage 4
 REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left,
 REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right,
 REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right,
 -- Stage 5
 REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right,
 REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right,
 -- Stage 6
 -- Stage 7
 REG_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 8
 REG_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 9
 REG_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 10
 REG_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 11
 REG_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 12
 REG_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 13
 REG_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 14
 REG_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 15
 REG_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 16
 REG_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 17
 REG_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 18
 REG_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 19
 REG_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 20
 REG_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 21
 REG_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 22
 REG_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 23
 REG_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 24
 REG_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 25
 REG_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 26
 REG_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 27
 REG_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 28
 REG_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 29
 REG_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 30
 REG_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 31
 REG_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 32
 REG_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 33
 REG_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 34
 REG_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 35
 REG_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 36
 REG_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 37
 REG_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 38
 REG_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 39
 REG_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 40
 REG_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 41
 REG_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 42
 REG_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 43
 REG_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 44
 REG_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 45
 REG_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 46
 REG_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 47
 REG_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 48
 REG_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 49
 REG_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 50
 REG_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 51
 REG_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 52
 REG_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 53
 REG_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 54
 REG_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 55
 REG_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 56
 REG_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 57
 REG_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 58
 REG_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 59
 REG_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 60
 REG_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 61
 REG_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 62
 REG_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 63
 REG_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 64
 REG_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 65
 REG_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 66
 REG_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 67
 REG_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 68
 REG_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 69
 REG_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 70
 REG_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 71
 REG_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 72
 REG_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 73
 REG_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 74
 REG_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 75
 REG_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 76
 REG_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 77
 REG_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 78
 REG_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 79
 REG_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 80
 REG_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 81
 REG_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 82
 REG_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 83
 REG_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 84
 REG_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 85
 REG_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 86
 REG_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 87
 REG_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 88
 REG_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 89
 REG_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 90
 REG_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 91
 REG_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 92
 REG_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 93
 REG_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 94
 REG_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 95
 REG_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 96
 REG_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 97
 REG_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 98
 REG_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 99
 REG_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 100
 REG_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 101
 REG_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 102
 REG_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 103
 REG_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 104
 REG_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 105
 REG_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 106
 REG_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 107
 REG_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 108
 REG_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 109
 REG_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 110
 REG_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 111
 REG_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 112
 REG_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 113
 REG_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 114
 REG_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 115
 REG_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 116
 REG_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 117
 REG_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 118
 REG_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 119
 REG_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 120
 REG_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 121
 REG_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 122
 REG_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 123
 REG_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 124
 REG_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 125
 REG_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 126
 REG_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 127
 REG_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 128
 REG_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 129
 REG_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 130
 REG_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 131
 REG_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 132
 REG_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 133
 REG_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 134
 REG_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 135
 REG_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 136
 REG_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 137
 REG_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 138
 REG_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 139
 REG_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 140
 REG_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 141
 REG_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 142
 REG_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 143
 REG_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 144
 REG_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 145
 REG_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 146
 REG_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 147
 REG_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 148
 REG_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 149
 REG_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 150
 REG_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 151
 REG_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 152
 REG_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 153
 REG_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 154
 REG_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 155
 REG_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 156
 REG_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 157
 REG_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 158
 REG_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 159
 REG_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 160
 REG_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 161
 REG_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 162
 REG_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 163
 REG_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 164
 REG_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 165
 REG_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 166
 REG_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 167
 REG_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 168
 REG_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 169
 REG_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 170
 REG_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 171
 REG_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 172
 REG_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 173
 REG_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 174
 REG_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 175
 REG_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 176
 REG_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 177
 REG_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 178
 REG_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 179
 REG_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 180
 REG_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 181
 REG_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 182
 REG_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 183
 REG_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 184
 REG_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 185
 REG_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 186
 REG_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 187
 REG_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 188
 REG_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 189
 REG_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 190
 REG_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 191
 REG_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 192
 REG_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 193
 REG_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 194
 REG_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 195
 REG_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 196
 REG_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 197
 REG_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 198
 REG_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 199
 REG_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 200
 REG_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 201
 REG_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 202
 REG_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 203
 REG_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 204
 REG_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 205
 REG_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 206
 REG_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 207
 REG_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 208
 REG_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 209
 REG_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 210
 REG_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 211
 REG_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 212
 REG_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 213
 REG_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 214
 REG_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 215
 REG_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 216
 REG_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 217
 REG_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 218
 REG_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 219
 REG_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 220
 REG_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 221
 REG_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 222
 REG_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 223
 REG_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 224
 REG_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 225
 REG_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 226
 REG_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 227
 REG_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 228
 REG_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 229
 REG_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 230
 REG_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 231
 REG_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 232
 REG_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 233
 REG_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 234
 REG_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 235
 REG_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 236
 REG_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 237
 REG_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 238
 REG_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 239
 REG_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 240
 REG_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 241
 REG_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 242
 REG_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 243
 REG_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 244
 REG_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 245
 REG_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 246
 REG_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 247
 REG_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 248
 REG_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 249
 REG_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 250
 REG_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 251
 REG_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 252
 REG_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 253
 REG_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 254
 REG_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 255
 REG_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 256
 REG_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 257
 REG_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 258
 REG_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 259
 REG_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 260
 REG_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 261
 REG_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 262
 REG_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 263
 REG_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 264
 REG_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 265
 REG_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 266
 REG_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 267
 REG_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 268
 REG_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 269
 REG_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 270
 REG_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 271
 REG_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 272
 REG_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 273
 REG_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 274
 REG_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 275
 REG_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 276
 REG_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 277
 REG_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 278
 REG_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 279
 REG_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 280
 REG_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 281
 REG_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 282
 REG_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 283
 REG_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 284
 REG_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 285
 REG_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 286
 REG_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 287
 REG_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 288
 REG_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 289
 REG_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 290
 REG_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 291
 REG_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 292
 REG_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 293
 REG_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 294
 REG_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 295
 REG_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 296
 REG_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 297
 REG_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 298
 REG_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 299
 REG_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 300
 REG_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 301
 REG_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 302
 REG_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 303
 REG_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 304
 REG_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 305
 REG_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 306
 REG_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 307
 REG_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 308
 REG_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 309
 REG_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 310
 REG_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 311
 REG_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 312
 REG_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 313
 REG_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 314
 REG_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 315
 REG_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 316
 REG_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 317
 REG_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 318
 REG_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 319
 REG_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 320
 REG_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 321
 REG_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 322
 REG_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 323
 REG_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 324
 REG_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 325
 REG_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 326
 REG_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 327
 REG_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 328
 REG_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 329
 REG_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 330
 REG_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 331
 REG_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 332
 REG_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 333
 REG_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 334
 REG_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 335
 REG_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 336
 REG_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 337
 REG_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 338
 REG_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 339
 REG_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 340
 REG_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 341
 REG_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 342
 REG_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 343
 REG_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 344
 REG_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 345
 REG_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 346
 REG_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 347
 REG_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 348
 REG_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 349
 REG_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 350
 REG_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 351
 REG_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 352
 REG_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 353
 REG_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 354
 REG_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 355
 REG_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 356
 REG_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 357
 REG_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 358
 REG_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 359
 REG_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 360
 REG_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 361
 REG_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 362
 REG_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 363
 REG_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 364
 REG_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 365
 REG_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 -- Stage 366
 REG_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond,
 REG_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse,
 REG_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse,
 REG_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse,
 -- Stage 367
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output,
 BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output,
 CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output,
 BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output,
 fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output,
 fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output,
 fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output,
 fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output,
 fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output,
 fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output,
 fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output,
 fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output,
 BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output,
 CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output,
 BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output,
 BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output,
 BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output,
 BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output,
 BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output,
 BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output,
 BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output,
 BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output,
 BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output,
 BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output,
 BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output,
 BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output,
 BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output,
 BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output,
 pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output,
 pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output,
 pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output,
 render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output,
 CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output,
 CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output,
 CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output,
 BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output,
 MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output,
 BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output,
 MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output,
 BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output,
 MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : pixel_t;
 variable VAR_i : unsigned(15 downto 0);
 variable VAR_j : unsigned(15 downto 0);
 variable VAR_state : full_state_t;
 variable VAR_scene : scene_t;
 variable VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l529_c19_e293_return_output : scene_t;
 variable VAR_cx : signed(15 downto 0);
 variable VAR_CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output : signed(15 downto 0);
 variable VAR_CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_x : signed(15 downto 0);
 variable VAR_cx_tr_pipelinec_gen_c_l531_c3_20d8 : signed(15 downto 0);
 variable VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_left : signed(15 downto 0);
 variable VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_right : signed(12 downto 0);
 variable VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output : signed(16 downto 0);
 variable VAR_cy : signed(15 downto 0);
 variable VAR_CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output : signed(15 downto 0);
 variable VAR_CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_x : signed(15 downto 0);
 variable VAR_cy_tr_pipelinec_gen_c_l533_c3_e577 : signed(15 downto 0);
 variable VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_left : signed(12 downto 0);
 variable VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_right : signed(15 downto 0);
 variable VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output : signed(16 downto 0);
 variable VAR_W : std_logic_vector(22 downto 0);
 variable VAR_H : std_logic_vector(22 downto 0);
 variable VAR_x : fixed;
 variable VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_left : fixed;
 variable VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_right : fixed;
 variable VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_a : fixed;
 variable VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_shift : signed(5 downto 0);
 variable VAR_fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_a : signed(15 downto 0);
 variable VAR_fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output : fixed;
 variable VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output : fixed;
 variable VAR_fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_a : std_logic_vector(22 downto 0);
 variable VAR_fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output : fixed;
 variable VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output : fixed;
 variable VAR_y : fixed;
 variable VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_left : fixed;
 variable VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_right : fixed;
 variable VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_a : fixed;
 variable VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_shift : signed(5 downto 0);
 variable VAR_fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_a : signed(15 downto 0);
 variable VAR_fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output : fixed;
 variable VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output : fixed;
 variable VAR_fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_a : std_logic_vector(22 downto 0);
 variable VAR_fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output : fixed;
 variable VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output : fixed;
 variable VAR_pix : pixel_t;
 variable VAR_scorebar : unsigned(15 downto 0);
 variable VAR_scorebar_tr_pipelinec_gen_c_l542_c12_3da9_0 : unsigned(15 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_left : unsigned(22 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_scene_t_scorebar_d41d_tr_pipelinec_gen_c_l542_c58_167d_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output : unsigned(38 downto 0);
 variable VAR_CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output : unsigned(38 downto 0);
 variable VAR_CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_x : unsigned(38 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_right : unsigned(16 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_right : unsigned(5 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output : unsigned(0 downto 0);
 variable VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue : unsigned(7 downto 0);
 variable VAR_pix_b_tr_pipelinec_gen_c_l547_c5_f9c7 : unsigned(7 downto 0);
 variable VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse : unsigned(7 downto 0);
 variable VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output : unsigned(7 downto 0);
 variable VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
 variable VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue : unsigned(7 downto 0);
 variable VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse : unsigned(7 downto 0);
 variable VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output : unsigned(7 downto 0);
 variable VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
 variable VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue : unsigned(7 downto 0);
 variable VAR_pix_r_tr_pipelinec_gen_c_l545_c5_1475 : unsigned(7 downto 0);
 variable VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse : unsigned(7 downto 0);
 variable VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output : unsigned(7 downto 0);
 variable VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond : unsigned(0 downto 0);
 variable VAR_c : fixed3;
 variable VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_x : fixed;
 variable VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_y : fixed;
 variable VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output : fixed3;
 variable VAR_r : unsigned(15 downto 0);
 variable VAR_r_tr_pipelinec_gen_c_l551_c14_5ae3_0 : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int22_t_fixed3_x_f_d41d_tr_pipelinec_gen_c_l551_c20_cba9_return_output : signed(21 downto 0);
 variable VAR_CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output : signed(21 downto 0);
 variable VAR_CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_x : signed(21 downto 0);
 variable VAR_g : unsigned(15 downto 0);
 variable VAR_g_tr_pipelinec_gen_c_l552_c14_3a9c_0 : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int22_t_fixed3_y_f_d41d_tr_pipelinec_gen_c_l552_c20_0a76_return_output : signed(21 downto 0);
 variable VAR_CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output : signed(21 downto 0);
 variable VAR_CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_x : signed(21 downto 0);
 variable VAR_b : unsigned(15 downto 0);
 variable VAR_b_tr_pipelinec_gen_c_l553_c14_f5bb_0 : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int22_t_fixed3_z_f_d41d_tr_pipelinec_gen_c_l553_c20_d145_return_output : signed(21 downto 0);
 variable VAR_CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output : signed(21 downto 0);
 variable VAR_CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_x : signed(21 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_cond : unsigned(0 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_right : unsigned(8 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output : unsigned(0 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output : unsigned(7 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_cond : unsigned(0 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_right : unsigned(8 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output : unsigned(0 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output : unsigned(7 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_cond : unsigned(0 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_right : unsigned(8 downto 0);
 variable VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_pixel_t_pixel_t_787c_tr_pipelinec_gen_c_l558_c10_7874_return_output : pixel_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_right := resize(to_unsigned(20, 5), 6);
     VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iftrue := to_unsigned(255, 8);
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_right := to_unsigned(256, 9);
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_right := to_unsigned(0, 1);
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_right := to_unsigned(0, 1);
     VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_left := signed(std_logic_vector(resize(to_unsigned(1081, 11), 13)));
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_right := to_unsigned(0, 1);
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_right := to_unsigned(0, 1);
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_right := to_unsigned(0, 1);
     VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iftrue := to_unsigned(255, 8);
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue := to_unsigned(200, 8);
     VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_right := signed(std_logic_vector(resize(to_unsigned(1921, 11), 13)));
     VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iftrue := to_unsigned(255, 8);
     VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_left := resize(to_unsigned(259, 9), 23);
     VAR_fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_a := resize_float_e_m_t(to_slv(to_float(0.9481481481481481, 8, 23)),8,23,8,14);
     VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_shift := signed(std_logic_vector(resize(to_unsigned(11, 4), 6)));
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_right := to_unsigned(0, 1);
     VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_right := to_unsigned(10, 4);
     VAR_pix_b_tr_pipelinec_gen_c_l547_c5_f9c7 := resize(to_unsigned(0, 1), 8);
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue := VAR_pix_b_tr_pipelinec_gen_c_l547_c5_f9c7;
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_right := to_unsigned(256, 9);
     VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_left := to_unsigned(10, 4);
     VAR_pix_r_tr_pipelinec_gen_c_l545_c5_1475 := resize(to_unsigned(0, 1), 8);
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue := VAR_pix_r_tr_pipelinec_gen_c_l545_c5_1475;
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_right := to_unsigned(256, 9);
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_right := to_unsigned(10, 4);
     VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_shift := signed(std_logic_vector(resize(to_unsigned(11, 4), 6)));
     VAR_fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_a := resize_float_e_m_t(to_slv(to_float(0.9481481481481482, 8, 23)),8,23,8,14);
     -- fixed_make_from_double[tr_pipelinec_gen_c_l539_c70_69e8] LATENCY=0
     -- Inputs
     fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_a <= VAR_fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_a;
     -- Outputs
     VAR_fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output := fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output;

     -- fixed_make_from_double[tr_pipelinec_gen_c_l538_c70_46cc] LATENCY=0
     -- Inputs
     fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_a <= VAR_fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_a;
     -- Outputs
     VAR_fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output := fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output;

     -- Submodule level 1
     VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_right := VAR_fixed_make_from_double_tr_pipelinec_gen_c_l539_c70_69e8_return_output;
     VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_right := VAR_fixed_make_from_double_tr_pipelinec_gen_c_l538_c70_46cc_return_output;
 -- Reads from global variables
     VAR_state := global_to_module.state;
     -- Submodule level 0
     -- CONST_REF_RD_scene_t_full_state_t_scene_d41d[tr_pipelinec_gen_c_l529_c19_e293] LATENCY=0
     VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l529_c19_e293_return_output := VAR_state.scene;

     -- Submodule level 1
     -- CONST_REF_RD_uint16_t_scene_t_scorebar_d41d[tr_pipelinec_gen_c_l542_c58_167d] LATENCY=0
     VAR_CONST_REF_RD_uint16_t_scene_t_scorebar_d41d_tr_pipelinec_gen_c_l542_c58_167d_return_output := VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l529_c19_e293_return_output.scorebar;

     -- Submodule level 2
     VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_right := VAR_CONST_REF_RD_uint16_t_scene_t_scorebar_d41d_tr_pipelinec_gen_c_l542_c58_167d_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_i := i;
     VAR_j := j;

     -- Submodule level 0
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_left := VAR_i;
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left := VAR_i;
     VAR_CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_x := signed(std_logic_vector(resize(VAR_i, 16)));
     VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_left := VAR_j;
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_left := VAR_j;
     VAR_CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_x := signed(std_logic_vector(resize(VAR_j, 16)));
     -- BIN_OP_INFERRED_MULT[tr_pipelinec_gen_c_l542_c24_cc3d] LATENCY=2
     -- Inputs
     BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_left <= VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_left;
     BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_right <= VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_right;

     -- BIN_OP_LT[tr_pipelinec_gen_c_l544_c82_eedf] LATENCY=1
     -- Inputs
     BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_left <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_left;
     BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_right <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_right;

     -- CONST_SL_1[tr_pipelinec_gen_c_l532_c16_046d] LATENCY=0
     -- Inputs
     CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_x <= VAR_CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_x;
     -- Outputs
     VAR_CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output := CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output;

     -- CONST_SL_1[tr_pipelinec_gen_c_l530_c16_86ea] LATENCY=0
     -- Inputs
     CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_x <= VAR_CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_x;
     -- Outputs
     VAR_CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output := CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output;

     -- BIN_OP_GTE[tr_pipelinec_gen_c_l544_c12_1c23] LATENCY=1
     -- Inputs
     BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_left <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_left;
     BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_right <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_right;

     -- BIN_OP_GT[tr_pipelinec_gen_c_l544_c61_d9c5] LATENCY=1
     -- Inputs
     BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_left <= VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_left;
     BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_right <= VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_right;

     -- Submodule level 1
     VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_left := VAR_CONST_SL_1_tr_pipelinec_gen_c_l530_c16_86ea_return_output;
     VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_right := VAR_CONST_SL_1_tr_pipelinec_gen_c_l532_c16_046d_return_output;
     -- BIN_OP_MINUS[tr_pipelinec_gen_c_l531_c8_94ad] LATENCY=1
     -- Inputs
     BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_left <= VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_left;
     BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_right <= VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_right;

     -- BIN_OP_MINUS[tr_pipelinec_gen_c_l533_c9_4b79] LATENCY=1
     -- Inputs
     BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_left <= VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_left;
     BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_right <= VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_right;

     -- Write to comb signals
     COMB_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left := REG_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     -- Submodule outputs
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output := BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output;
     VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output := BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output;
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output := BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output;
     VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output := BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output;
     VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output := BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output;

     -- Submodule level 0
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_left := VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l544_c12_1c23_return_output;
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_left := VAR_BIN_OP_GT_tr_pipelinec_gen_c_l544_c61_d9c5_return_output;
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_left := VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c82_eedf_return_output;
     VAR_cx_tr_pipelinec_gen_c_l531_c3_20d8 := resize(VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l531_c8_94ad_return_output, 16);
     VAR_cy_tr_pipelinec_gen_c_l533_c3_e577 := resize(VAR_BIN_OP_MINUS_tr_pipelinec_gen_c_l533_c9_4b79_return_output, 16);
     VAR_fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_a := VAR_cx_tr_pipelinec_gen_c_l531_c3_20d8;
     VAR_fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_a := VAR_cy_tr_pipelinec_gen_c_l533_c3_e577;
     -- fixed_make_from_short[tr_pipelinec_gen_c_l538_c33_b52e] LATENCY=0
     -- Inputs
     fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_a <= VAR_fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_a;
     -- Outputs
     VAR_fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output := fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output;

     -- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c82_478a] LATENCY=0
     -- Inputs
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_left <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_left;
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_right <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_right;
     -- Outputs
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output := BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output;

     -- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c12_5895] LATENCY=0
     -- Inputs
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_left <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_left;
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_right <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_right;
     -- Outputs
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output := BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output;

     -- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c61_beb7] LATENCY=0
     -- Inputs
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_left <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_left;
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_right <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_right;
     -- Outputs
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output := BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output;

     -- fixed_make_from_short[tr_pipelinec_gen_c_l539_c33_31d5] LATENCY=0
     -- Inputs
     fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_a <= VAR_fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_a;
     -- Outputs
     VAR_fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output := fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output;

     -- Submodule level 1
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left := VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_5895_return_output;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right := VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c61_beb7_return_output;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right := VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c82_478a_return_output;
     VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_a := VAR_fixed_make_from_short_tr_pipelinec_gen_c_l538_c33_b52e_return_output;
     VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_a := VAR_fixed_make_from_short_tr_pipelinec_gen_c_l539_c33_31d5_return_output;
     -- fixed_shr[tr_pipelinec_gen_c_l539_c23_7550] LATENCY=0
     -- Inputs
     fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_a <= VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_a;
     fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_shift <= VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_shift;
     -- Outputs
     VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output := fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output;

     -- fixed_shr[tr_pipelinec_gen_c_l538_c23_82ce] LATENCY=0
     -- Inputs
     fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_a <= VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_a;
     fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_shift <= VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_shift;
     -- Outputs
     VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output := fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output;

     -- Submodule level 2
     VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_left := VAR_fixed_shr_tr_pipelinec_gen_c_l538_c23_82ce_return_output;
     VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_left := VAR_fixed_shr_tr_pipelinec_gen_c_l539_c23_7550_return_output;
     -- fixed_mul[tr_pipelinec_gen_c_l539_c13_9a90] LATENCY=5
     -- Inputs
     fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_left <= VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_left;
     fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_right <= VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_right;

     -- fixed_mul[tr_pipelinec_gen_c_l538_c13_ffb3] LATENCY=5
     -- Inputs
     fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_left <= VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_left;
     fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_right <= VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_right;

     -- Write to comb signals
     COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     COMB_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left := REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left := REG_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right := REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right := REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Submodule outputs
     VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output := BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output;

     -- Submodule level 0
     VAR_CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_x := VAR_BIN_OP_INFERRED_MULT_tr_pipelinec_gen_c_l542_c24_cc3d_return_output;
     -- CONST_SR_11[tr_pipelinec_gen_c_l542_c24_cb53] LATENCY=0
     -- Inputs
     CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_x <= VAR_CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_x;
     -- Outputs
     VAR_CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output := CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output;

     -- Submodule level 1
     VAR_scorebar_tr_pipelinec_gen_c_l542_c12_3da9_0 := resize(VAR_CONST_SR_11_tr_pipelinec_gen_c_l542_c24_cb53_return_output, 16);
     VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_right := VAR_scorebar_tr_pipelinec_gen_c_l542_c12_3da9_0;
     -- BIN_OP_PLUS[tr_pipelinec_gen_c_l544_c33_633d] LATENCY=1
     -- Inputs
     BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_left <= VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_left;
     BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_right <= VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_right;

     -- Write to comb signals
     COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     COMB_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left := REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left := REG_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right := REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right := REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Submodule outputs
     VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output := BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output;

     -- Submodule level 0
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_right := VAR_BIN_OP_PLUS_tr_pipelinec_gen_c_l544_c33_633d_return_output;
     -- BIN_OP_LT[tr_pipelinec_gen_c_l544_c29_d00f] LATENCY=1
     -- Inputs
     BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_right <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_right;

     -- Write to comb signals
     COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left := REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right := REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right := REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Submodule outputs
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output := BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output;

     -- Submodule level 0
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_left := VAR_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_return_output;
     -- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c29_766f] LATENCY=1
     -- Inputs
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_left <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_left;
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_right <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_right;

     -- Write to comb signals
     COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left := REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right := REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right := REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Submodule outputs
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output := BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output;

     -- Submodule level 0
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_right := VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c29_766f_return_output;
     -- BIN_OP_AND[tr_pipelinec_gen_c_l544_c12_48d6] LATENCY=0
     -- Inputs
     BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_right;
     -- Outputs
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output := BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output;

     -- Submodule level 1
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_left := VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_return_output;
     -- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c12_ae4d] LATENCY=1
     -- Inputs
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_left <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_left;
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_right <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_right;

     -- Write to comb signals
     COMB_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     COMB_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right := REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right := REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Submodule outputs
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output := BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output;
     VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output := fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output;
     VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output := fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output;

     -- Submodule level 0
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_left := VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_ae4d_return_output;
     VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_x := VAR_fixed_mul_tr_pipelinec_gen_c_l538_c13_ffb3_return_output;
     VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_y := VAR_fixed_mul_tr_pipelinec_gen_c_l539_c13_9a90_return_output;
     -- BIN_OP_AND[tr_pipelinec_gen_c_l544_c12_925a] LATENCY=0
     -- Inputs
     BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_left;
     BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     -- Outputs
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output := BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output;

     -- render_pixel_internal[tr_pipelinec_gen_c_l550_c16_85da] LATENCY=360
     -- Inputs
     render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_x <= VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_x;
     render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_y <= VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_y;

     -- Submodule level 1
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_left := VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_return_output;
     -- BIN_OP_NEQ[tr_pipelinec_gen_c_l544_c12_6cb4] LATENCY=0
     -- Inputs
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_left <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_left;
     BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_right <= VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_right;
     -- Outputs
     VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output := BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output;

     -- Submodule level 2
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_left := VAR_BIN_OP_NEQ_tr_pipelinec_gen_c_l544_c12_6cb4_return_output;
     -- BIN_OP_AND[tr_pipelinec_gen_c_l544_c12_d8f8] LATENCY=1
     -- Inputs
     BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_left <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_left;
     BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;

     -- Write to comb signals
   elsif STAGE = 7 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output := BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output;

     -- Submodule level 0
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := VAR_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_return_output;
     -- Write to comb signals
     COMB_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 13 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 14 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 15 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 16 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 17 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 18 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 19 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 20 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 21 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 22 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 23 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 24 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 25 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 26 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 27 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 28 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 29 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 30 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 31 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 32 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 33 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 34 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 35 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 36 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 37 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 38 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 39 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 40 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 41 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 42 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 43 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 44 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 45 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 46 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 47 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 48 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 49 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 50 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 51 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 52 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 53 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 54 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 55 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 56 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 57 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 58 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 59 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 60 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 61 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 62 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 63 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 64 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 65 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 66 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 67 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 68 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 69 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 70 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 71 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 72 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 73 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 74 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 75 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 76 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 77 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 78 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 79 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 80 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 81 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 82 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 83 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 84 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 85 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 86 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 87 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 88 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 89 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 90 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 91 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 92 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 93 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 94 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 95 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 96 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 97 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 98 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 99 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 100 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 101 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 102 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 103 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 104 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 105 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 106 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 107 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 108 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 109 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 110 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 111 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 112 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 113 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 114 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 115 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 116 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 117 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 118 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 119 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 120 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 121 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 122 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 123 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 124 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 125 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 126 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 127 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 128 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 129 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 130 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 131 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 132 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 133 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 134 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 135 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 136 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 137 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 138 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 139 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 140 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 141 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 142 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 143 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 144 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 145 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 146 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 147 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 148 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 149 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 150 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 151 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 152 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 153 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 154 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 155 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 156 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 157 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 158 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 159 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 160 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 161 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 162 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 163 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 164 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 165 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 166 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 167 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 168 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 169 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 170 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 171 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 172 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 173 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 174 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 175 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 176 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 177 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 178 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 179 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 180 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 181 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 182 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 183 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 184 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 185 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 186 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 187 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 188 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 189 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 190 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 191 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 192 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 193 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 194 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 195 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 196 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 197 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 198 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 199 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 200 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 201 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 202 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 203 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 204 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 205 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 206 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 207 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 208 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 209 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 210 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 211 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 212 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 213 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 214 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 215 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 216 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 217 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 218 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 219 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 220 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 221 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 222 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 223 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 224 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 225 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 226 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 227 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 228 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 229 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 230 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 231 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 232 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 233 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 234 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 235 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 236 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 237 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 238 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 239 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 240 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 241 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 242 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 243 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 244 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 245 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 246 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 247 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 248 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 249 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 250 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 251 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 252 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 253 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 254 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 255 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 256 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 257 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 258 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 259 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 260 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 261 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 262 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 263 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 264 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 265 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 266 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 267 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 268 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 269 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 270 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 271 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 272 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 273 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 274 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 275 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 276 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 277 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 278 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 279 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 280 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 281 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 282 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 283 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 284 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 285 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 286 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 287 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 288 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 289 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 290 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 291 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 292 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 293 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 294 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 295 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 296 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 297 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 298 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 299 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 300 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 301 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 302 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 303 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 304 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 305 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 306 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 307 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 308 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 309 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 310 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 311 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 312 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 313 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 314 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 315 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 316 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 317 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 318 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 319 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 320 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 321 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 322 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 323 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 324 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 325 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 326 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 327 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 328 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 329 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 330 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 331 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 332 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 333 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 334 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 335 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 336 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 337 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 338 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 339 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 340 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 341 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 342 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 343 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 344 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 345 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 346 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 347 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 348 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 349 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 350 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 351 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 352 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 353 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 354 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 355 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 356 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 357 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 358 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 359 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 360 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 361 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 362 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 363 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 364 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 365 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;

     -- Write to comb signals
     COMB_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
   elsif STAGE = 366 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Submodule outputs
     VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output := render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_int22_t_fixed3_y_f_d41d[tr_pipelinec_gen_c_l552_c20_0a76] LATENCY=0
     VAR_CONST_REF_RD_int22_t_fixed3_y_f_d41d_tr_pipelinec_gen_c_l552_c20_0a76_return_output := VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output.y.f;

     -- CONST_REF_RD_int22_t_fixed3_z_f_d41d[tr_pipelinec_gen_c_l553_c20_d145] LATENCY=0
     VAR_CONST_REF_RD_int22_t_fixed3_z_f_d41d_tr_pipelinec_gen_c_l553_c20_d145_return_output := VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output.z.f;

     -- CONST_REF_RD_int22_t_fixed3_x_f_d41d[tr_pipelinec_gen_c_l551_c20_cba9] LATENCY=0
     VAR_CONST_REF_RD_int22_t_fixed3_x_f_d41d_tr_pipelinec_gen_c_l551_c20_cba9_return_output := VAR_render_pixel_internal_tr_pipelinec_gen_c_l550_c16_85da_return_output.x.f;

     -- Submodule level 1
     VAR_CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_x := VAR_CONST_REF_RD_int22_t_fixed3_x_f_d41d_tr_pipelinec_gen_c_l551_c20_cba9_return_output;
     VAR_CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_x := VAR_CONST_REF_RD_int22_t_fixed3_y_f_d41d_tr_pipelinec_gen_c_l552_c20_0a76_return_output;
     VAR_CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_x := VAR_CONST_REF_RD_int22_t_fixed3_z_f_d41d_tr_pipelinec_gen_c_l553_c20_d145_return_output;
     -- CONST_SR_2[tr_pipelinec_gen_c_l551_c20_29b3] LATENCY=0
     -- Inputs
     CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_x <= VAR_CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_x;
     -- Outputs
     VAR_CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output := CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output;

     -- CONST_SR_2[tr_pipelinec_gen_c_l553_c20_6ab8] LATENCY=0
     -- Inputs
     CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_x <= VAR_CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_x;
     -- Outputs
     VAR_CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output := CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output;

     -- CONST_SR_2[tr_pipelinec_gen_c_l552_c20_c1b4] LATENCY=0
     -- Inputs
     CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_x <= VAR_CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_x;
     -- Outputs
     VAR_CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output := CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output;

     -- Submodule level 2
     VAR_r_tr_pipelinec_gen_c_l551_c14_5ae3_0 := resize(unsigned(std_logic_vector(VAR_CONST_SR_2_tr_pipelinec_gen_c_l551_c20_29b3_return_output)),16);
     VAR_g_tr_pipelinec_gen_c_l552_c14_3a9c_0 := resize(unsigned(std_logic_vector(VAR_CONST_SR_2_tr_pipelinec_gen_c_l552_c20_c1b4_return_output)),16);
     VAR_b_tr_pipelinec_gen_c_l553_c14_f5bb_0 := resize(unsigned(std_logic_vector(VAR_CONST_SR_2_tr_pipelinec_gen_c_l553_c20_6ab8_return_output)),16);
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_left := VAR_b_tr_pipelinec_gen_c_l553_c14_f5bb_0;
     VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse := resize(VAR_b_tr_pipelinec_gen_c_l553_c14_f5bb_0, 8);
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_left := VAR_g_tr_pipelinec_gen_c_l552_c14_3a9c_0;
     VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse := resize(VAR_g_tr_pipelinec_gen_c_l552_c14_3a9c_0, 8);
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_left := VAR_r_tr_pipelinec_gen_c_l551_c14_5ae3_0;
     VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse := resize(VAR_r_tr_pipelinec_gen_c_l551_c14_5ae3_0, 8);
     -- BIN_OP_GTE[tr_pipelinec_gen_c_l554_c14_8e81] LATENCY=1
     -- Inputs
     BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_left <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_left;
     BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_right <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_right;

     -- BIN_OP_GTE[tr_pipelinec_gen_c_l556_c14_374a] LATENCY=1
     -- Inputs
     BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_left <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_left;
     BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_right <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_right;

     -- BIN_OP_GTE[tr_pipelinec_gen_c_l555_c14_77f4] LATENCY=1
     -- Inputs
     BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_left <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_left;
     BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_right <= VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_right;

     -- Write to comb signals
     COMB_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     COMB_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse <= VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse;
     COMB_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse <= VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse;
     COMB_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse <= VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse;
   elsif STAGE = 367 then
     -- Read from prev stage
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond := REG_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse := REG_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse;
     VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse := REG_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse;
     VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse := REG_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse;
     -- Submodule outputs
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output := BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output;
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output := BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output;
     VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output := BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output;

     -- Submodule level 0
     VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_cond := VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l554_c14_8e81_return_output;
     VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_cond := VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l555_c14_77f4_return_output;
     VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_cond := VAR_BIN_OP_GTE_tr_pipelinec_gen_c_l556_c14_374a_return_output;
     -- MUX[tr_pipelinec_gen_c_l555_c14_6d28] LATENCY=0
     -- Inputs
     MUX_tr_pipelinec_gen_c_l555_c14_6d28_cond <= VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_cond;
     MUX_tr_pipelinec_gen_c_l555_c14_6d28_iftrue <= VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iftrue;
     MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse <= VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse;
     -- Outputs
     VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output := MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output;

     -- MUX[tr_pipelinec_gen_c_l556_c14_02b9] LATENCY=0
     -- Inputs
     MUX_tr_pipelinec_gen_c_l556_c14_02b9_cond <= VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_cond;
     MUX_tr_pipelinec_gen_c_l556_c14_02b9_iftrue <= VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iftrue;
     MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse <= VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse;
     -- Outputs
     VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output := MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output;

     -- MUX[tr_pipelinec_gen_c_l554_c14_f66a] LATENCY=0
     -- Inputs
     MUX_tr_pipelinec_gen_c_l554_c14_f66a_cond <= VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_cond;
     MUX_tr_pipelinec_gen_c_l554_c14_f66a_iftrue <= VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iftrue;
     MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse <= VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse;
     -- Outputs
     VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output := MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output;

     -- Submodule level 1
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse := VAR_MUX_tr_pipelinec_gen_c_l554_c14_f66a_return_output;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse := VAR_MUX_tr_pipelinec_gen_c_l555_c14_6d28_return_output;
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse := VAR_MUX_tr_pipelinec_gen_c_l556_c14_02b9_return_output;
     -- pix_b_MUX[tr_pipelinec_gen_c_l544_c3_e881] LATENCY=1
     -- Inputs
     pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue;
     pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse <= VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse;

     -- pix_g_MUX[tr_pipelinec_gen_c_l544_c3_e881] LATENCY=1
     -- Inputs
     pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue;
     pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse <= VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse;

     -- pix_r_MUX[tr_pipelinec_gen_c_l544_c3_e881] LATENCY=1
     -- Inputs
     pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iftrue;
     pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse <= VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_iffalse;

     -- Write to comb signals
   elsif STAGE = 368 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output := pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output;
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output := pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output;
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output := pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_pixel_t_pixel_t_787c[tr_pipelinec_gen_c_l558_c10_7874] LATENCY=0
     VAR_CONST_REF_RD_pixel_t_pixel_t_787c_tr_pipelinec_gen_c_l558_c10_7874_return_output := CONST_REF_RD_pixel_t_pixel_t_787c(
     pixel_t_NULL,
     VAR_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output,
     VAR_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output,
     VAR_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_return_output);

     -- Submodule level 1
     VAR_return_output := VAR_CONST_REF_RD_pixel_t_pixel_t_787c_tr_pipelinec_gen_c_l558_c10_7874_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= COMB_STAGE0_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     -- Stage 1
     REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     REG_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= COMB_STAGE1_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     REG_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= COMB_STAGE1_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Stage 2
     REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     REG_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left <= COMB_STAGE2_BIN_OP_LT_tr_pipelinec_gen_c_l544_c29_d00f_left;
     REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     REG_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= COMB_STAGE2_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Stage 3
     REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     REG_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= COMB_STAGE3_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Stage 4
     REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left <= COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_48d6_left;
     REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     REG_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= COMB_STAGE4_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Stage 5
     REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right <= COMB_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_925a_right;
     REG_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right <= COMB_STAGE5_BIN_OP_AND_tr_pipelinec_gen_c_l544_c12_d8f8_right;
     -- Stage 6
     -- Stage 7
     REG_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE7_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE7_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE7_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 8
     REG_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE8_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE8_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE8_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 9
     REG_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE9_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE9_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE9_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 10
     REG_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE10_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE10_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE10_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 11
     REG_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE11_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE11_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE11_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 12
     REG_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE12_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE12_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE12_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 13
     REG_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE13_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE13_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE13_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 14
     REG_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE14_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE14_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE14_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 15
     REG_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE15_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE15_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE15_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 16
     REG_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE16_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE16_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE16_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 17
     REG_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE17_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE17_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE17_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 18
     REG_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE18_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE18_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE18_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 19
     REG_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE19_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE19_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE19_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 20
     REG_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE20_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE20_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE20_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 21
     REG_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE21_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE21_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE21_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 22
     REG_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE22_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE22_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE22_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 23
     REG_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE23_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE23_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE23_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 24
     REG_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE24_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE24_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE24_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 25
     REG_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE25_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE25_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE25_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 26
     REG_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE26_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE26_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE26_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 27
     REG_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE27_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE27_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE27_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 28
     REG_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE28_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE28_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE28_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 29
     REG_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE29_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE29_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE29_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 30
     REG_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE30_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE30_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE30_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 31
     REG_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE31_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE31_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE31_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 32
     REG_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE32_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE32_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE32_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 33
     REG_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE33_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE33_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE33_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 34
     REG_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE34_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE34_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE34_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 35
     REG_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE35_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE35_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE35_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 36
     REG_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE36_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE36_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE36_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 37
     REG_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE37_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE37_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE37_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 38
     REG_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE38_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE38_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE38_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 39
     REG_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE39_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE39_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE39_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 40
     REG_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE40_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE40_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE40_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 41
     REG_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE41_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE41_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE41_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 42
     REG_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE42_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE42_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE42_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 43
     REG_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE43_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE43_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE43_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 44
     REG_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE44_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE44_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE44_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 45
     REG_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE45_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE45_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE45_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 46
     REG_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE46_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE46_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE46_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 47
     REG_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE47_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE47_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE47_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 48
     REG_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE48_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE48_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE48_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 49
     REG_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE49_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE49_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE49_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 50
     REG_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE50_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE50_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE50_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 51
     REG_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE51_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE51_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE51_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 52
     REG_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE52_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE52_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE52_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 53
     REG_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE53_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE53_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE53_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 54
     REG_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE54_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE54_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE54_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 55
     REG_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE55_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE55_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE55_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 56
     REG_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE56_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE56_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE56_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 57
     REG_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE57_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE57_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE57_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 58
     REG_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE58_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE58_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE58_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 59
     REG_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE59_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE59_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE59_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 60
     REG_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE60_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE60_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE60_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 61
     REG_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE61_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE61_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE61_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 62
     REG_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE62_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE62_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE62_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 63
     REG_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE63_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE63_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE63_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 64
     REG_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE64_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE64_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE64_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 65
     REG_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE65_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE65_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE65_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 66
     REG_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE66_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE66_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE66_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 67
     REG_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE67_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE67_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE67_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 68
     REG_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE68_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE68_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE68_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 69
     REG_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE69_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE69_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE69_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 70
     REG_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE70_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE70_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE70_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 71
     REG_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE71_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE71_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE71_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 72
     REG_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE72_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE72_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE72_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 73
     REG_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE73_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE73_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE73_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 74
     REG_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE74_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE74_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE74_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 75
     REG_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE75_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE75_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE75_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 76
     REG_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE76_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE76_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE76_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 77
     REG_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE77_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE77_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE77_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 78
     REG_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE78_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE78_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE78_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 79
     REG_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE79_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE79_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE79_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 80
     REG_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE80_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE80_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE80_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 81
     REG_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE81_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE81_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE81_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 82
     REG_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE82_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE82_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE82_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 83
     REG_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE83_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE83_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE83_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 84
     REG_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE84_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE84_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE84_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 85
     REG_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE85_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE85_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE85_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 86
     REG_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE86_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE86_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE86_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 87
     REG_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE87_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE87_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE87_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 88
     REG_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE88_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE88_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE88_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 89
     REG_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE89_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE89_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE89_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 90
     REG_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE90_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE90_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE90_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 91
     REG_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE91_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE91_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE91_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 92
     REG_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE92_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE92_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE92_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 93
     REG_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE93_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE93_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE93_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 94
     REG_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE94_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE94_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE94_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 95
     REG_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE95_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE95_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE95_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 96
     REG_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE96_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE96_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE96_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 97
     REG_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE97_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE97_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE97_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 98
     REG_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE98_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE98_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE98_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 99
     REG_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE99_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE99_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE99_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 100
     REG_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE100_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE100_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE100_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 101
     REG_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE101_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE101_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE101_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 102
     REG_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE102_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE102_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE102_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 103
     REG_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE103_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE103_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE103_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 104
     REG_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE104_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE104_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE104_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 105
     REG_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE105_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE105_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE105_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 106
     REG_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE106_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE106_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE106_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 107
     REG_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE107_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE107_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE107_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 108
     REG_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE108_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE108_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE108_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 109
     REG_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE109_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE109_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE109_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 110
     REG_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE110_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE110_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE110_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 111
     REG_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE111_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE111_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE111_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 112
     REG_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE112_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE112_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE112_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 113
     REG_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE113_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE113_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE113_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 114
     REG_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE114_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE114_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE114_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 115
     REG_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE115_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE115_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE115_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 116
     REG_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE116_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE116_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE116_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 117
     REG_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE117_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE117_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE117_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 118
     REG_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE118_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE118_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE118_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 119
     REG_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE119_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE119_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE119_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 120
     REG_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE120_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE120_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE120_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 121
     REG_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE121_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE121_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE121_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 122
     REG_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE122_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE122_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE122_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 123
     REG_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE123_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE123_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE123_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 124
     REG_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE124_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE124_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE124_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 125
     REG_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE125_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE125_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE125_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 126
     REG_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE126_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE126_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE126_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 127
     REG_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE127_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE127_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE127_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 128
     REG_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE128_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE128_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE128_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 129
     REG_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE129_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE129_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE129_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 130
     REG_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE130_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE130_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE130_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 131
     REG_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE131_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE131_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE131_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 132
     REG_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE132_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE132_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE132_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 133
     REG_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE133_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE133_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE133_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 134
     REG_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE134_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE134_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE134_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 135
     REG_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE135_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE135_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE135_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 136
     REG_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE136_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE136_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE136_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 137
     REG_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE137_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE137_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE137_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 138
     REG_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE138_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE138_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE138_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 139
     REG_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE139_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE139_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE139_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 140
     REG_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE140_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE140_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE140_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 141
     REG_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE141_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE141_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE141_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 142
     REG_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE142_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE142_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE142_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 143
     REG_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE143_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE143_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE143_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 144
     REG_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE144_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE144_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE144_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 145
     REG_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE145_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE145_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE145_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 146
     REG_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE146_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE146_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE146_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 147
     REG_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE147_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE147_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE147_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 148
     REG_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE148_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE148_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE148_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 149
     REG_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE149_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE149_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE149_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 150
     REG_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE150_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE150_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE150_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 151
     REG_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE151_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE151_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE151_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 152
     REG_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE152_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE152_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE152_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 153
     REG_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE153_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE153_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE153_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 154
     REG_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE154_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE154_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE154_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 155
     REG_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE155_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE155_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE155_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 156
     REG_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE156_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE156_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE156_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 157
     REG_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE157_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE157_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE157_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 158
     REG_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE158_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE158_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE158_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 159
     REG_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE159_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE159_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE159_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 160
     REG_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE160_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE160_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE160_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 161
     REG_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE161_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE161_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE161_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 162
     REG_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE162_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE162_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE162_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 163
     REG_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE163_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE163_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE163_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 164
     REG_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE164_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE164_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE164_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 165
     REG_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE165_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE165_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE165_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 166
     REG_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE166_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE166_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE166_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 167
     REG_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE167_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE167_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE167_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 168
     REG_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE168_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE168_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE168_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 169
     REG_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE169_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE169_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE169_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 170
     REG_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE170_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE170_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE170_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 171
     REG_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE171_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE171_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE171_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 172
     REG_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE172_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE172_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE172_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 173
     REG_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE173_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE173_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE173_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 174
     REG_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE174_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE174_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE174_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 175
     REG_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE175_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE175_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE175_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 176
     REG_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE176_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE176_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE176_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 177
     REG_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE177_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE177_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE177_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 178
     REG_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE178_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE178_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE178_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 179
     REG_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE179_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE179_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE179_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 180
     REG_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE180_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE180_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE180_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 181
     REG_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE181_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE181_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE181_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 182
     REG_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE182_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE182_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE182_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 183
     REG_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE183_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE183_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE183_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 184
     REG_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE184_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE184_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE184_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 185
     REG_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE185_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE185_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE185_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 186
     REG_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE186_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE186_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE186_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 187
     REG_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE187_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE187_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE187_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 188
     REG_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE188_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE188_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE188_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 189
     REG_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE189_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE189_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE189_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 190
     REG_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE190_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE190_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE190_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 191
     REG_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE191_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE191_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE191_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 192
     REG_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE192_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE192_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE192_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 193
     REG_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE193_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE193_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE193_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 194
     REG_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE194_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE194_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE194_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 195
     REG_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE195_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE195_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE195_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 196
     REG_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE196_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE196_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE196_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 197
     REG_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE197_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE197_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE197_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 198
     REG_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE198_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE198_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE198_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 199
     REG_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE199_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE199_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE199_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 200
     REG_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE200_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE200_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE200_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 201
     REG_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE201_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE201_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE201_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 202
     REG_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE202_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE202_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE202_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 203
     REG_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE203_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE203_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE203_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 204
     REG_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE204_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE204_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE204_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 205
     REG_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE205_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE205_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE205_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 206
     REG_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE206_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE206_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE206_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 207
     REG_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE207_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE207_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE207_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 208
     REG_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE208_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE208_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE208_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 209
     REG_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE209_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE209_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE209_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 210
     REG_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE210_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE210_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE210_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 211
     REG_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE211_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE211_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE211_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 212
     REG_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE212_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE212_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE212_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 213
     REG_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE213_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE213_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE213_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 214
     REG_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE214_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE214_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE214_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 215
     REG_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE215_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE215_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE215_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 216
     REG_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE216_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE216_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE216_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 217
     REG_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE217_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE217_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE217_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 218
     REG_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE218_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE218_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE218_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 219
     REG_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE219_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE219_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE219_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 220
     REG_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE220_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE220_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE220_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 221
     REG_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE221_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE221_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE221_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 222
     REG_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE222_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE222_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE222_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 223
     REG_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE223_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE223_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE223_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 224
     REG_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE224_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE224_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE224_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 225
     REG_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE225_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE225_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE225_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 226
     REG_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE226_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE226_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE226_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 227
     REG_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE227_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE227_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE227_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 228
     REG_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE228_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE228_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE228_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 229
     REG_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE229_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE229_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE229_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 230
     REG_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE230_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE230_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE230_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 231
     REG_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE231_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE231_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE231_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 232
     REG_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE232_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE232_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE232_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 233
     REG_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE233_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE233_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE233_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 234
     REG_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE234_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE234_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE234_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 235
     REG_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE235_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE235_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE235_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 236
     REG_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE236_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE236_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE236_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 237
     REG_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE237_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE237_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE237_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 238
     REG_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE238_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE238_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE238_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 239
     REG_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE239_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE239_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE239_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 240
     REG_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE240_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE240_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE240_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 241
     REG_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE241_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE241_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE241_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 242
     REG_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE242_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE242_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE242_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 243
     REG_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE243_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE243_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE243_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 244
     REG_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE244_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE244_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE244_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 245
     REG_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE245_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE245_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE245_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 246
     REG_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE246_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE246_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE246_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 247
     REG_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE247_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE247_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE247_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 248
     REG_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE248_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE248_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE248_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 249
     REG_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE249_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE249_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE249_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 250
     REG_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE250_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE250_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE250_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 251
     REG_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE251_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE251_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE251_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 252
     REG_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE252_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE252_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE252_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 253
     REG_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE253_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE253_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE253_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 254
     REG_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE254_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE254_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE254_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 255
     REG_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE255_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE255_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE255_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 256
     REG_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE256_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE256_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE256_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 257
     REG_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE257_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE257_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE257_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 258
     REG_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE258_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE258_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE258_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 259
     REG_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE259_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE259_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE259_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 260
     REG_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE260_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE260_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE260_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 261
     REG_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE261_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE261_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE261_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 262
     REG_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE262_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE262_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE262_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 263
     REG_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE263_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE263_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE263_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 264
     REG_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE264_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE264_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE264_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 265
     REG_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE265_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE265_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE265_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 266
     REG_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE266_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE266_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE266_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 267
     REG_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE267_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE267_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE267_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 268
     REG_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE268_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE268_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE268_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 269
     REG_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE269_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE269_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE269_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 270
     REG_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE270_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE270_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE270_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 271
     REG_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE271_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE271_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE271_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 272
     REG_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE272_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE272_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE272_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 273
     REG_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE273_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE273_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE273_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 274
     REG_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE274_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE274_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE274_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 275
     REG_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE275_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE275_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE275_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 276
     REG_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE276_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE276_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE276_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 277
     REG_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE277_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE277_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE277_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 278
     REG_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE278_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE278_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE278_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 279
     REG_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE279_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE279_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE279_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 280
     REG_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE280_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE280_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE280_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 281
     REG_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE281_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE281_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE281_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 282
     REG_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE282_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE282_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE282_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 283
     REG_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE283_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE283_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE283_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 284
     REG_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE284_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE284_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE284_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 285
     REG_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE285_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE285_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE285_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 286
     REG_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE286_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE286_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE286_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 287
     REG_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE287_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE287_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE287_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 288
     REG_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE288_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE288_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE288_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 289
     REG_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE289_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE289_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE289_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 290
     REG_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE290_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE290_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE290_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 291
     REG_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE291_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE291_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE291_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 292
     REG_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE292_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE292_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE292_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 293
     REG_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE293_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE293_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE293_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 294
     REG_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE294_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE294_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE294_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 295
     REG_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE295_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE295_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE295_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 296
     REG_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE296_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE296_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE296_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 297
     REG_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE297_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE297_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE297_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 298
     REG_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE298_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE298_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE298_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 299
     REG_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE299_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE299_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE299_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 300
     REG_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE300_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE300_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE300_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 301
     REG_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE301_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE301_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE301_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 302
     REG_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE302_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE302_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE302_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 303
     REG_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE303_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE303_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE303_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 304
     REG_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE304_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE304_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE304_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 305
     REG_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE305_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE305_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE305_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 306
     REG_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE306_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE306_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE306_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 307
     REG_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE307_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE307_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE307_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 308
     REG_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE308_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE308_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE308_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 309
     REG_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE309_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE309_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE309_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 310
     REG_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE310_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE310_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE310_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 311
     REG_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE311_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE311_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE311_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 312
     REG_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE312_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE312_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE312_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 313
     REG_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE313_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE313_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE313_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 314
     REG_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE314_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE314_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE314_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 315
     REG_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE315_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE315_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE315_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 316
     REG_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE316_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE316_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE316_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 317
     REG_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE317_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE317_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE317_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 318
     REG_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE318_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE318_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE318_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 319
     REG_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE319_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE319_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE319_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 320
     REG_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE320_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE320_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE320_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 321
     REG_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE321_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE321_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE321_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 322
     REG_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE322_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE322_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE322_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 323
     REG_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE323_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE323_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE323_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 324
     REG_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE324_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE324_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE324_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 325
     REG_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE325_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE325_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE325_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 326
     REG_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE326_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE326_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE326_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 327
     REG_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE327_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE327_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE327_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 328
     REG_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE328_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE328_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE328_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 329
     REG_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE329_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE329_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE329_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 330
     REG_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE330_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE330_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE330_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 331
     REG_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE331_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE331_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE331_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 332
     REG_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE332_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE332_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE332_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 333
     REG_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE333_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE333_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE333_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 334
     REG_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE334_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE334_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE334_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 335
     REG_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE335_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE335_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE335_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 336
     REG_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE336_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE336_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE336_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 337
     REG_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE337_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE337_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE337_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 338
     REG_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE338_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE338_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE338_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 339
     REG_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE339_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE339_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE339_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 340
     REG_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE340_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE340_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE340_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 341
     REG_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE341_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE341_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE341_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 342
     REG_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE342_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE342_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE342_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 343
     REG_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE343_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE343_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE343_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 344
     REG_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE344_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE344_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE344_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 345
     REG_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE345_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE345_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE345_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 346
     REG_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE346_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE346_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE346_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 347
     REG_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE347_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE347_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE347_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 348
     REG_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE348_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE348_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE348_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 349
     REG_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE349_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE349_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE349_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 350
     REG_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE350_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE350_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE350_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 351
     REG_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE351_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE351_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE351_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 352
     REG_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE352_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE352_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE352_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 353
     REG_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE353_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE353_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE353_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 354
     REG_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE354_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE354_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE354_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 355
     REG_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE355_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE355_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE355_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 356
     REG_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE356_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE356_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE356_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 357
     REG_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE357_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE357_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE357_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 358
     REG_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE358_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE358_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE358_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 359
     REG_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE359_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE359_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE359_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 360
     REG_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE360_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE360_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE360_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 361
     REG_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE361_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE361_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE361_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 362
     REG_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE362_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE362_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE362_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 363
     REG_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE363_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE363_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE363_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 364
     REG_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE364_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE364_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE364_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 365
     REG_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE365_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE365_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE365_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     -- Stage 366
     REG_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE366_pix_b_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE366_pix_g_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond <= COMB_STAGE366_pix_r_MUX_tr_pipelinec_gen_c_l544_c3_e881_cond;
     REG_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse <= COMB_STAGE366_MUX_tr_pipelinec_gen_c_l554_c14_f66a_iffalse;
     REG_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse <= COMB_STAGE366_MUX_tr_pipelinec_gen_c_l555_c14_6d28_iffalse;
     REG_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse <= COMB_STAGE366_MUX_tr_pipelinec_gen_c_l556_c14_02b9_iffalse;
     -- Stage 367
 end if;
end process;

end arch;
