-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.003453985168853315, 0.007939485626724333, 0.012424986084595356, 0.01691048654246637, 0.02139598700033739, 0.025881487458208414, 0.030366987916079433, 0.03485248837395044, 0.039337988831821456, 0.04382348928969248, 0.048308989747563494, 0.05279449020543452, 0.057279990663305545, 0.061765491121176574, 0.0662509915790476, 0.07073649203691862, 0.07522199249478964, 0.07970749295266068, 0.0841929934105317, 0.08867849386840272, 0.09316399432627373, 0.09764949478414477, 0.1021349952420158, 0.10662049569988684, 0.11110599615775783, 0.11559149661562884, 0.12007699707349985, 0.12456249753137086, 0.12904799798924185, 0.1335334984471129, 0.1380189989049839, 0.14250449936285492, 0.14698999982072594, 0.15147550027859696, 0.15596100073646793, 0.16044650119433895, 0.16493200165220995, 0.16941750211008097, 0.17390300256795196, 0.178388503025823, 0.18287400348369398, 0.187359503941565, 0.191845004399436, 0.19633050485730702, 0.20081600531517807, 0.20530150577304906, 0.2097870062309201, 0.21427250668879108, 0.2187580071466621, 0.2232435076045331, 0.22772900806240412, 0.23221450852027511, 0.23670000897814616, 0.24118550943601721, 0.24567100989388826, 0.2501565103517593, 0.2546420108096303, 0.25912751126750133, 0.2636130117253724, 0.26809851218324343, 0.2725840126411145, 0.27706951309898553, 0.2815550135568566, 0.2860405140147276, 0.29052601447259857, 0.2950115149304697, 0.2994970153883407, 0.3039825158462118, 0.3084680163040828, 0.3129535167619539, 0.31743901721982487, 0.321924517677696, 0.32641001813556697, 0.33089551859343797, 0.33538101905130896, 0.33986651950918, 0.34435201996705106, 0.34883752042492205, 0.35332302088279316, 0.35780852134066427, 0.36229402179853526, 0.3667795222564063, 0.37126502271427736, 0.3757505231721484, 0.3802360236300194, 0.38472152408789045, 0.3892070245457615, 0.39369252500363255, 0.39817802546150355, 0.40266352591937454, 0.40714902637724565, 0.41163452683511664, 0.41612002729298764, 0.4206055277508588, 0.4250910282087298, 0.42957652866660084, 0.4340620291244719, 0.4385475295823429, 0.443033030040214, 0.447518530498085, 0.4520040309559561, 0.4564895314138271, 0.4609750318716981, 0.46546053232956913, 0.4699460327874401, 0.4744315332453112, 0.4789170337031823, 0.4834025341610533, 0.4878880346189244, 0.4923735350767954, 0.49685903553466637, 0.5013445359925374, 0.5058300364504084, 0.5103155369082794, 0.5148010373661502, 0.5192865378240212, 0.5237720382818923, 0.5282575387397632, 0.5327430391976342, 0.5372285396555052, 0.5417140401133762, 0.5461995405712472, 0.5506850410291181, 0.5551705414869892, 0.5596560419448602, 0.5641415424027311, 0.5686270428606021, 0.5731125433184731, 0.577598043776344, 0.582083544234215, 0.586569044692086, 0.591054545149957, 0.595540045607828, 0.6000255460656989, 0.6045110465235699, 0.6089965469814409, 0.6134820474393119, 0.6179675478971829, 0.6224530483550539, 0.6269385488129249, 0.6314240492707959, 0.6359095497286668, 0.6403950501865378, 0.6448805506444089, 0.6493660511022799, 0.6538515515601508, 0.6583370520180217, 0.6628225524758925, 0.6673080529337636, 0.6717935533916346, 0.6762790538495057, 0.6807645543073766, 0.6852500547652476, 0.6897355552231186, 0.6942210556809896, 0.6987065561388606, 0.7031920565967315, 0.7076775570546024, 0.7121630575124736, 0.7166485579703443, 0.7211340584282153, 0.7256195588860864, 0.7301050593439574, 0.7345905598018284, 0.7390760602596994, 0.7435615607175704, 0.7480470611754414, 0.7525325616333123, 0.7570180620911833, 0.7615035625490543, 0.7659890630069253, 0.7704745634647964, 0.7749600639226671, 0.7794455643805382, 0.783931064838409, 0.78841656529628, 0.7929020657541511, 0.7973875662120222, 0.8018730666698931, 0.8063585671277641, 0.8108440675856351, 0.8153295680435061, 0.8198150685013771, 0.8243005689592481, 0.828786069417119, 0.8332715698749898, 0.8377570703328608, 0.8422425707907318, 0.8467280712486029, 0.8512135717064739, 0.8556990721643447, 0.8601845726222159, 0.8646700730800869, 0.8691555735379579, 0.8736410739958289, 0.8781265744536998, 0.8826120749115708, 0.8870975753694418, 0.8915830758273127, 0.8960685762851837, 0.9005540767430547, 0.9050395772009255, 0.9095250776587965, 0.9140105781166675, 0.9184960785745387, 0.9229815790324096, 0.9274670794902806, 0.9319525799481516, 0.9364380804060226, 0.9409235808638936, 0.9454090813217646, 0.9498945817796355, 0.9543800822375064, 0.9588655826953774, 0.9633510831532484, 0.9678365836111193, 0.9723220840689905, 0.9768075845268614, 0.9812930849847324, 0.9857785854426034, 0.9902640859004744, 0.9947495863583454, 0.9992350868162163]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 7
entity render_pixel_internal_360CLK_987815b4 is
port(
 clk : in std_logic;
 global_to_module : in render_pixel_internal_global_to_module_t;
 x : in fixed;
 y : in fixed;
 return_output : out fixed3);
end render_pixel_internal_360CLK_987815b4;
architecture arch of render_pixel_internal_360CLK_987815b4 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 360;
-- All of the wires/regs in function
-- Stage 0
-- Stage 1
-- Stage 2
-- Stage 3
signal REG_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 4
signal REG_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 5
signal REG_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 6
signal REG_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 7
signal REG_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 8
signal REG_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 9
signal REG_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 10
signal REG_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 11
signal REG_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 12
signal REG_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 13
signal REG_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 14
signal REG_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 15
signal REG_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 16
signal REG_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 17
signal REG_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 18
signal REG_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 19
signal REG_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 20
signal REG_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 21
signal REG_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 22
signal REG_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 23
signal REG_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 24
signal REG_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 25
signal REG_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 26
signal REG_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 27
signal REG_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 28
signal REG_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 29
signal REG_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 30
signal REG_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 31
signal REG_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 32
signal REG_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 33
signal REG_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 34
signal REG_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 35
signal REG_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 36
signal REG_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
signal COMB_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
-- Stage 37
-- Stage 38
-- Stage 39
-- Stage 40
-- Stage 41
-- Stage 42
-- Stage 43
-- Stage 44
-- Stage 45
-- Stage 46
-- Stage 47
-- Stage 48
-- Stage 49
-- Stage 50
-- Stage 51
-- Stage 52
-- Stage 53
-- Stage 54
-- Stage 55
-- Stage 56
-- Stage 57
-- Stage 58
-- Stage 59
-- Stage 60
-- Stage 61
-- Stage 62
-- Stage 63
-- Stage 64
-- Stage 65
-- Stage 66
-- Stage 67
-- Stage 68
-- Stage 69
-- Stage 70
-- Stage 71
-- Stage 72
-- Stage 73
-- Stage 74
-- Stage 75
-- Stage 76
-- Stage 77
-- Stage 78
-- Stage 79
-- Stage 80
-- Stage 81
-- Stage 82
-- Stage 83
-- Stage 84
-- Stage 85
-- Stage 86
-- Stage 87
-- Stage 88
-- Stage 89
-- Stage 90
-- Stage 91
-- Stage 92
-- Stage 93
-- Stage 94
-- Stage 95
-- Stage 96
-- Stage 97
-- Stage 98
-- Stage 99
-- Stage 100
-- Stage 101
-- Stage 102
-- Stage 103
-- Stage 104
-- Stage 105
-- Stage 106
-- Stage 107
-- Stage 108
-- Stage 109
-- Stage 110
-- Stage 111
-- Stage 112
-- Stage 113
-- Stage 114
-- Stage 115
-- Stage 116
-- Stage 117
-- Stage 118
-- Stage 119
-- Stage 120
-- Stage 121
-- Stage 122
-- Stage 123
-- Stage 124
-- Stage 125
-- Stage 126
-- Stage 127
-- Stage 128
-- Stage 129
-- Stage 130
-- Stage 131
-- Stage 132
-- Stage 133
-- Stage 134
-- Stage 135
-- Stage 136
-- Stage 137
-- Stage 138
-- Stage 139
-- Stage 140
-- Stage 141
-- Stage 142
-- Stage 143
-- Stage 144
-- Stage 145
-- Stage 146
-- Stage 147
-- Stage 148
-- Stage 149
-- Stage 150
-- Stage 151
-- Stage 152
-- Stage 153
-- Stage 154
-- Stage 155
-- Stage 156
-- Stage 157
-- Stage 158
-- Stage 159
-- Stage 160
-- Stage 161
-- Stage 162
-- Stage 163
-- Stage 164
-- Stage 165
-- Stage 166
-- Stage 167
-- Stage 168
-- Stage 169
-- Stage 170
-- Stage 171
-- Stage 172
-- Stage 173
-- Stage 174
-- Stage 175
-- Stage 176
-- Stage 177
-- Stage 178
-- Stage 179
-- Stage 180
-- Stage 181
-- Stage 182
-- Stage 183
-- Stage 184
-- Stage 185
-- Stage 186
-- Stage 187
-- Stage 188
-- Stage 189
-- Stage 190
-- Stage 191
-- Stage 192
-- Stage 193
-- Stage 194
-- Stage 195
-- Stage 196
-- Stage 197
-- Stage 198
-- Stage 199
-- Stage 200
-- Stage 201
-- Stage 202
-- Stage 203
-- Stage 204
-- Stage 205
-- Stage 206
-- Stage 207
-- Stage 208
-- Stage 209
-- Stage 210
-- Stage 211
-- Stage 212
-- Stage 213
-- Stage 214
-- Stage 215
-- Stage 216
-- Stage 217
-- Stage 218
-- Stage 219
-- Stage 220
-- Stage 221
-- Stage 222
-- Stage 223
-- Stage 224
-- Stage 225
-- Stage 226
-- Stage 227
-- Stage 228
-- Stage 229
-- Stage 230
-- Stage 231
-- Stage 232
-- Stage 233
-- Stage 234
-- Stage 235
-- Stage 236
-- Stage 237
-- Stage 238
-- Stage 239
-- Stage 240
-- Stage 241
-- Stage 242
-- Stage 243
-- Stage 244
-- Stage 245
-- Stage 246
-- Stage 247
-- Stage 248
-- Stage 249
-- Stage 250
-- Stage 251
-- Stage 252
-- Stage 253
-- Stage 254
-- Stage 255
-- Stage 256
-- Stage 257
-- Stage 258
-- Stage 259
-- Stage 260
-- Stage 261
-- Stage 262
-- Stage 263
-- Stage 264
-- Stage 265
-- Stage 266
-- Stage 267
-- Stage 268
-- Stage 269
-- Stage 270
-- Stage 271
-- Stage 272
-- Stage 273
-- Stage 274
-- Stage 275
-- Stage 276
-- Stage 277
-- Stage 278
-- Stage 279
-- Stage 280
-- Stage 281
-- Stage 282
-- Stage 283
-- Stage 284
-- Stage 285
-- Stage 286
-- Stage 287
-- Stage 288
-- Stage 289
-- Stage 290
-- Stage 291
-- Stage 292
-- Stage 293
-- Stage 294
-- Stage 295
-- Stage 296
-- Stage 297
-- Stage 298
-- Stage 299
-- Stage 300
-- Stage 301
-- Stage 302
-- Stage 303
-- Stage 304
-- Stage 305
-- Stage 306
-- Stage 307
-- Stage 308
-- Stage 309
-- Stage 310
-- Stage 311
-- Stage 312
-- Stage 313
-- Stage 314
-- Stage 315
-- Stage 316
-- Stage 317
-- Stage 318
-- Stage 319
-- Stage 320
-- Stage 321
-- Stage 322
-- Stage 323
-- Stage 324
-- Stage 325
-- Stage 326
-- Stage 327
-- Stage 328
-- Stage 329
-- Stage 330
-- Stage 331
-- Stage 332
-- Stage 333
-- Stage 334
-- Stage 335
-- Stage 336
-- Stage 337
-- Stage 338
-- Stage 339
-- Stage 340
-- Stage 341
-- Stage 342
-- Stage 343
-- Stage 344
-- Stage 345
-- Stage 346
-- Stage 347
-- Stage 348
-- Stage 349
-- Stage 350
-- Stage 351
-- Stage 352
-- Stage 353
-- Stage 354
-- Stage 355
-- Stage 356
-- Stage 357
-- Stage 358
-- Stage 359
-- Each function instance gets signals
-- object_coord_to_float3[tr_pipelinec_gen_c_l422_c16_ccf5]
signal object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_a : fixed3;
signal object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;

-- fixed_to_float[tr_pipelinec_gen_c_l423_c24_ab0b]
signal fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_a : fixed;
signal fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output : std_logic_vector(22 downto 0);

-- fixed_to_float[tr_pipelinec_gen_c_l423_c43_dd5f]
signal fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_a : fixed;
signal fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output : std_logic_vector(22 downto 0);

-- normalize[tr_pipelinec_gen_c_l424_c15_c26c]
signal normalize_tr_pipelinec_gen_c_l424_c15_c26c_v : float3;
signal normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output : float3;

-- cast_ray[tr_pipelinec_gen_c_l425_c10_8f9f]
signal cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_hitin : point_and_dir;
signal cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output : fixed3;

function CONST_REF_RD_float3_float3_7d4c( ref_toks_0 : std_logic_vector;
 ref_toks_1 : std_logic_vector;
 ref_toks_2 : std_logic_vector) return float3 is
 
  variable base : float3; 
  variable return_output : float3;
begin
      base.x := ref_toks_0;
      base.y := ref_toks_1;
      base.z := ref_toks_2;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_point_and_dir_point_and_dir_8057( ref_toks_0 : float3;
 ref_toks_1 : float3) return point_and_dir is
 
  variable base : point_and_dir; 
  variable return_output : point_and_dir;
begin
      base.orig := ref_toks_0;
      base.dir := ref_toks_1;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5
object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5 : entity work.object_coord_to_float3_3CLK_9d26212c port map (
clk,
object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_a,
object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output);

-- fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b
fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b : entity work.fixed_to_float_3CLK_adafa2ea port map (
clk,
fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_a,
fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output);

-- fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f
fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f : entity work.fixed_to_float_3CLK_adafa2ea port map (
clk,
fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_a,
fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output);

-- normalize_tr_pipelinec_gen_c_l424_c15_c26c
normalize_tr_pipelinec_gen_c_l424_c15_c26c : entity work.normalize_34CLK_495496ce port map (
clk,
normalize_tr_pipelinec_gen_c_l424_c15_c26c_v,
normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output);

-- cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f
cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f : entity work.cast_ray_323CLK_f2c1ab37 port map (
clk,
global_to_module.cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f,
cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_hitin,
cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 x,
 y,
 -- Registers
 -- Stage 0
 -- Stage 1
 -- Stage 2
 -- Stage 3
 REG_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 4
 REG_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 5
 REG_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 6
 REG_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 7
 REG_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 8
 REG_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 9
 REG_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 10
 REG_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 11
 REG_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 12
 REG_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 13
 REG_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 14
 REG_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 15
 REG_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 16
 REG_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 17
 REG_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 18
 REG_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 19
 REG_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 20
 REG_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 21
 REG_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 22
 REG_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 23
 REG_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 24
 REG_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 25
 REG_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 26
 REG_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 27
 REG_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 28
 REG_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 29
 REG_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 30
 REG_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 31
 REG_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 32
 REG_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 33
 REG_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 34
 REG_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 35
 REG_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 36
 REG_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 -- Stage 37
 -- Stage 38
 -- Stage 39
 -- Stage 40
 -- Stage 41
 -- Stage 42
 -- Stage 43
 -- Stage 44
 -- Stage 45
 -- Stage 46
 -- Stage 47
 -- Stage 48
 -- Stage 49
 -- Stage 50
 -- Stage 51
 -- Stage 52
 -- Stage 53
 -- Stage 54
 -- Stage 55
 -- Stage 56
 -- Stage 57
 -- Stage 58
 -- Stage 59
 -- Stage 60
 -- Stage 61
 -- Stage 62
 -- Stage 63
 -- Stage 64
 -- Stage 65
 -- Stage 66
 -- Stage 67
 -- Stage 68
 -- Stage 69
 -- Stage 70
 -- Stage 71
 -- Stage 72
 -- Stage 73
 -- Stage 74
 -- Stage 75
 -- Stage 76
 -- Stage 77
 -- Stage 78
 -- Stage 79
 -- Stage 80
 -- Stage 81
 -- Stage 82
 -- Stage 83
 -- Stage 84
 -- Stage 85
 -- Stage 86
 -- Stage 87
 -- Stage 88
 -- Stage 89
 -- Stage 90
 -- Stage 91
 -- Stage 92
 -- Stage 93
 -- Stage 94
 -- Stage 95
 -- Stage 96
 -- Stage 97
 -- Stage 98
 -- Stage 99
 -- Stage 100
 -- Stage 101
 -- Stage 102
 -- Stage 103
 -- Stage 104
 -- Stage 105
 -- Stage 106
 -- Stage 107
 -- Stage 108
 -- Stage 109
 -- Stage 110
 -- Stage 111
 -- Stage 112
 -- Stage 113
 -- Stage 114
 -- Stage 115
 -- Stage 116
 -- Stage 117
 -- Stage 118
 -- Stage 119
 -- Stage 120
 -- Stage 121
 -- Stage 122
 -- Stage 123
 -- Stage 124
 -- Stage 125
 -- Stage 126
 -- Stage 127
 -- Stage 128
 -- Stage 129
 -- Stage 130
 -- Stage 131
 -- Stage 132
 -- Stage 133
 -- Stage 134
 -- Stage 135
 -- Stage 136
 -- Stage 137
 -- Stage 138
 -- Stage 139
 -- Stage 140
 -- Stage 141
 -- Stage 142
 -- Stage 143
 -- Stage 144
 -- Stage 145
 -- Stage 146
 -- Stage 147
 -- Stage 148
 -- Stage 149
 -- Stage 150
 -- Stage 151
 -- Stage 152
 -- Stage 153
 -- Stage 154
 -- Stage 155
 -- Stage 156
 -- Stage 157
 -- Stage 158
 -- Stage 159
 -- Stage 160
 -- Stage 161
 -- Stage 162
 -- Stage 163
 -- Stage 164
 -- Stage 165
 -- Stage 166
 -- Stage 167
 -- Stage 168
 -- Stage 169
 -- Stage 170
 -- Stage 171
 -- Stage 172
 -- Stage 173
 -- Stage 174
 -- Stage 175
 -- Stage 176
 -- Stage 177
 -- Stage 178
 -- Stage 179
 -- Stage 180
 -- Stage 181
 -- Stage 182
 -- Stage 183
 -- Stage 184
 -- Stage 185
 -- Stage 186
 -- Stage 187
 -- Stage 188
 -- Stage 189
 -- Stage 190
 -- Stage 191
 -- Stage 192
 -- Stage 193
 -- Stage 194
 -- Stage 195
 -- Stage 196
 -- Stage 197
 -- Stage 198
 -- Stage 199
 -- Stage 200
 -- Stage 201
 -- Stage 202
 -- Stage 203
 -- Stage 204
 -- Stage 205
 -- Stage 206
 -- Stage 207
 -- Stage 208
 -- Stage 209
 -- Stage 210
 -- Stage 211
 -- Stage 212
 -- Stage 213
 -- Stage 214
 -- Stage 215
 -- Stage 216
 -- Stage 217
 -- Stage 218
 -- Stage 219
 -- Stage 220
 -- Stage 221
 -- Stage 222
 -- Stage 223
 -- Stage 224
 -- Stage 225
 -- Stage 226
 -- Stage 227
 -- Stage 228
 -- Stage 229
 -- Stage 230
 -- Stage 231
 -- Stage 232
 -- Stage 233
 -- Stage 234
 -- Stage 235
 -- Stage 236
 -- Stage 237
 -- Stage 238
 -- Stage 239
 -- Stage 240
 -- Stage 241
 -- Stage 242
 -- Stage 243
 -- Stage 244
 -- Stage 245
 -- Stage 246
 -- Stage 247
 -- Stage 248
 -- Stage 249
 -- Stage 250
 -- Stage 251
 -- Stage 252
 -- Stage 253
 -- Stage 254
 -- Stage 255
 -- Stage 256
 -- Stage 257
 -- Stage 258
 -- Stage 259
 -- Stage 260
 -- Stage 261
 -- Stage 262
 -- Stage 263
 -- Stage 264
 -- Stage 265
 -- Stage 266
 -- Stage 267
 -- Stage 268
 -- Stage 269
 -- Stage 270
 -- Stage 271
 -- Stage 272
 -- Stage 273
 -- Stage 274
 -- Stage 275
 -- Stage 276
 -- Stage 277
 -- Stage 278
 -- Stage 279
 -- Stage 280
 -- Stage 281
 -- Stage 282
 -- Stage 283
 -- Stage 284
 -- Stage 285
 -- Stage 286
 -- Stage 287
 -- Stage 288
 -- Stage 289
 -- Stage 290
 -- Stage 291
 -- Stage 292
 -- Stage 293
 -- Stage 294
 -- Stage 295
 -- Stage 296
 -- Stage 297
 -- Stage 298
 -- Stage 299
 -- Stage 300
 -- Stage 301
 -- Stage 302
 -- Stage 303
 -- Stage 304
 -- Stage 305
 -- Stage 306
 -- Stage 307
 -- Stage 308
 -- Stage 309
 -- Stage 310
 -- Stage 311
 -- Stage 312
 -- Stage 313
 -- Stage 314
 -- Stage 315
 -- Stage 316
 -- Stage 317
 -- Stage 318
 -- Stage 319
 -- Stage 320
 -- Stage 321
 -- Stage 322
 -- Stage 323
 -- Stage 324
 -- Stage 325
 -- Stage 326
 -- Stage 327
 -- Stage 328
 -- Stage 329
 -- Stage 330
 -- Stage 331
 -- Stage 332
 -- Stage 333
 -- Stage 334
 -- Stage 335
 -- Stage 336
 -- Stage 337
 -- Stage 338
 -- Stage 339
 -- Stage 340
 -- Stage 341
 -- Stage 342
 -- Stage 343
 -- Stage 344
 -- Stage 345
 -- Stage 346
 -- Stage 347
 -- Stage 348
 -- Stage 349
 -- Stage 350
 -- Stage 351
 -- Stage 352
 -- Stage 353
 -- Stage 354
 -- Stage 355
 -- Stage 356
 -- Stage 357
 -- Stage 358
 -- Stage 359
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
 fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output,
 fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output,
 normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output,
 cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : fixed3;
 variable VAR_x : fixed;
 variable VAR_y : fixed;
 variable VAR_state : full_state_t;
 variable VAR_scene : scene_t;
 variable VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l419_c19_0b43_return_output : scene_t;
 variable VAR_colors : scene_colors_t;
 variable VAR_hitin : point_and_dir;
 variable VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_a : fixed3;
 variable VAR_CONST_REF_RD_fixed3_scene_t_camera_d41d_tr_pipelinec_gen_c_l422_c39_a24f_return_output : fixed3;
 variable VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output : float3;
 variable VAR_camera_dir : float3;
 variable VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_a : fixed;
 variable VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output : std_logic_vector(22 downto 0);
 variable VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_a : fixed;
 variable VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output : std_logic_vector(22 downto 0);
 variable VAR_normalize_tr_pipelinec_gen_c_l424_c15_c26c_v : float3;
 variable VAR_CONST_REF_RD_float3_float3_7d4c_tr_pipelinec_gen_c_l424_c25_c910_return_output : float3;
 variable VAR_normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output : float3;
 variable VAR_cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_hitin : point_and_dir;
 variable VAR_CONST_REF_RD_point_and_dir_point_and_dir_8057_tr_pipelinec_gen_c_l425_c19_8a0d_return_output : point_and_dir;
 variable VAR_cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output : fixed3;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
 -- Reads from global variables
     VAR_state := global_to_module.state;
     -- Submodule level 0
     -- CONST_REF_RD_scene_t_full_state_t_scene_d41d[tr_pipelinec_gen_c_l419_c19_0b43] LATENCY=0
     VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l419_c19_0b43_return_output := VAR_state.scene;

     -- Submodule level 1
     -- CONST_REF_RD_fixed3_scene_t_camera_d41d[tr_pipelinec_gen_c_l422_c39_a24f] LATENCY=0
     VAR_CONST_REF_RD_fixed3_scene_t_camera_d41d_tr_pipelinec_gen_c_l422_c39_a24f_return_output := VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l419_c19_0b43_return_output.camera;

     -- Submodule level 2
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_a := VAR_CONST_REF_RD_fixed3_scene_t_camera_d41d_tr_pipelinec_gen_c_l422_c39_a24f_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_x := x;
     VAR_y := y;

     -- Submodule level 0
     VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_a := VAR_x;
     VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_a := VAR_y;
     -- object_coord_to_float3[tr_pipelinec_gen_c_l422_c16_ccf5] LATENCY=3
     -- Inputs
     object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_a <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_a;

     -- fixed_to_float[tr_pipelinec_gen_c_l423_c24_ab0b] LATENCY=3
     -- Inputs
     fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_a <= VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_a;

     -- fixed_to_float[tr_pipelinec_gen_c_l423_c43_dd5f] LATENCY=3
     -- Inputs
     fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_a <= VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_a;

     -- Write to comb signals
   elsif STAGE = 1 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 2 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 3 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output := fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output;
     VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output := fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output;
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_float3_float3_7d4c[tr_pipelinec_gen_c_l424_c25_c910] LATENCY=0
     VAR_CONST_REF_RD_float3_float3_7d4c_tr_pipelinec_gen_c_l424_c25_c910_return_output := CONST_REF_RD_float3_float3_7d4c(
     VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c24_ab0b_return_output,
     VAR_fixed_to_float_tr_pipelinec_gen_c_l423_c43_dd5f_return_output,
     to_slv(to_float(-1.0, 8, 14)));

     -- Submodule level 1
     VAR_normalize_tr_pipelinec_gen_c_l424_c15_c26c_v := VAR_CONST_REF_RD_float3_float3_7d4c_tr_pipelinec_gen_c_l424_c25_c910_return_output;
     -- normalize[tr_pipelinec_gen_c_l424_c15_c26c] LATENCY=34
     -- Inputs
     normalize_tr_pipelinec_gen_c_l424_c15_c26c_v <= VAR_normalize_tr_pipelinec_gen_c_l424_c15_c26c_v;

     -- Write to comb signals
     COMB_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 7 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 13 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 14 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 15 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 16 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 17 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 18 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 19 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 20 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 21 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 22 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 23 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 24 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 25 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 26 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 27 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 28 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 29 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 30 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 31 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 32 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 33 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 34 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 35 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 36 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;

     -- Write to comb signals
     COMB_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
   elsif STAGE = 37 then
     -- Read from prev stage
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output := REG_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Submodule outputs
     VAR_normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output := normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_point_and_dir_point_and_dir_8057[tr_pipelinec_gen_c_l425_c19_8a0d] LATENCY=0
     VAR_CONST_REF_RD_point_and_dir_point_and_dir_8057_tr_pipelinec_gen_c_l425_c19_8a0d_return_output := CONST_REF_RD_point_and_dir_point_and_dir_8057(
     VAR_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output,
     VAR_normalize_tr_pipelinec_gen_c_l424_c15_c26c_return_output);

     -- Submodule level 1
     VAR_cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_hitin := VAR_CONST_REF_RD_point_and_dir_point_and_dir_8057_tr_pipelinec_gen_c_l425_c19_8a0d_return_output;
     -- cast_ray[tr_pipelinec_gen_c_l425_c10_8f9f] LATENCY=323
     -- Inputs
     cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_hitin <= VAR_cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_hitin;

     -- Write to comb signals
   elsif STAGE = 38 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 39 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 40 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 41 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 42 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 43 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 44 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 45 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 46 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 47 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 48 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 49 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 50 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 51 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 52 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 53 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 54 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 55 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 56 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 57 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 58 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 59 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 60 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 61 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 62 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 63 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 64 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 65 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 66 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 67 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 68 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 69 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 70 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 71 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 72 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 73 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 74 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 75 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 76 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 77 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 78 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 79 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 80 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 81 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 82 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 83 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 84 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 85 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 86 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 87 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 88 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 89 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 90 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 91 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 92 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 93 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 94 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 95 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 96 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 97 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 98 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 99 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 100 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 101 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 102 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 103 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 104 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 105 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 106 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 107 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 108 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 109 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 110 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 111 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 112 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 113 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 114 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 115 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 116 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 117 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 118 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 119 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 120 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 121 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 122 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 123 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 124 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 125 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 126 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 127 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 128 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 129 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 130 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 131 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 132 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 133 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 134 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 135 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 136 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 137 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 138 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 139 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 140 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 141 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 142 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 143 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 144 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 145 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 146 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 147 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 148 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 149 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 150 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 151 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 152 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 153 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 154 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 155 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 156 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 157 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 158 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 159 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 160 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 161 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 162 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 163 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 164 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 165 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 166 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 167 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 168 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 169 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 170 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 171 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 172 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 173 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 174 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 175 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 176 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 177 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 178 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 179 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 180 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 181 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 182 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 183 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 184 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 185 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 186 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 187 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 188 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 189 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 190 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 191 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 192 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 193 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 194 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 195 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 196 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 197 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 198 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 199 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 200 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 201 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 202 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 203 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 204 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 205 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 206 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 207 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 208 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 209 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 210 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 211 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 212 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 213 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 214 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 215 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 216 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 217 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 218 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 219 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 220 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 221 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 222 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 223 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 224 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 225 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 226 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 227 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 228 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 229 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 230 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 231 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 232 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 233 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 234 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 235 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 236 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 237 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 238 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 239 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 240 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 241 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 242 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 243 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 244 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 245 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 246 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 247 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 248 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 249 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 250 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 251 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 252 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 253 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 254 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 255 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 256 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 257 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 258 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 259 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 260 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 261 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 262 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 263 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 264 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 265 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 266 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 267 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 268 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 269 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 270 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 271 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 272 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 273 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 274 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 275 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 276 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 277 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 278 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 279 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 280 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 281 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 282 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 283 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 284 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 285 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 286 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 287 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 288 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 289 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 290 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 291 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 292 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 293 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 294 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 295 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 296 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 297 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 298 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 299 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 300 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 301 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 302 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 303 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 304 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 305 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 306 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 307 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 308 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 309 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 310 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 311 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 312 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 313 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 314 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 315 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 316 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 317 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 318 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 319 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 320 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 321 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 322 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 323 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 324 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 325 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 326 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 327 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 328 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 329 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 330 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 331 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 332 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 333 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 334 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 335 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 336 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 337 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 338 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 339 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 340 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 341 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 342 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 343 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 344 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 345 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 346 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 347 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 348 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 349 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 350 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 351 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 352 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 353 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 354 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 355 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 356 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 357 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 358 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 359 then
     -- Read from prev stage

     -- Write to comb signals
   elsif STAGE = 360 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output := cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output;

     -- Submodule level 0
     VAR_return_output := VAR_cast_ray_tr_pipelinec_gen_c_l425_c10_8f9f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     -- Stage 1
     -- Stage 2
     -- Stage 3
     REG_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE3_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 4
     REG_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE4_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 5
     REG_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE5_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 6
     REG_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE6_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 7
     REG_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE7_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 8
     REG_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE8_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 9
     REG_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE9_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 10
     REG_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE10_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 11
     REG_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE11_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 12
     REG_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE12_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 13
     REG_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE13_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 14
     REG_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE14_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 15
     REG_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE15_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 16
     REG_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE16_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 17
     REG_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE17_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 18
     REG_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE18_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 19
     REG_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE19_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 20
     REG_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE20_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 21
     REG_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE21_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 22
     REG_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE22_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 23
     REG_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE23_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 24
     REG_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE24_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 25
     REG_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE25_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 26
     REG_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE26_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 27
     REG_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE27_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 28
     REG_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE28_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 29
     REG_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE29_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 30
     REG_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE30_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 31
     REG_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE31_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 32
     REG_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE32_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 33
     REG_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE33_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 34
     REG_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE34_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 35
     REG_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE35_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 36
     REG_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output <= COMB_STAGE36_object_coord_to_float3_tr_pipelinec_gen_c_l422_c16_ccf5_return_output;
     -- Stage 37
     -- Stage 38
     -- Stage 39
     -- Stage 40
     -- Stage 41
     -- Stage 42
     -- Stage 43
     -- Stage 44
     -- Stage 45
     -- Stage 46
     -- Stage 47
     -- Stage 48
     -- Stage 49
     -- Stage 50
     -- Stage 51
     -- Stage 52
     -- Stage 53
     -- Stage 54
     -- Stage 55
     -- Stage 56
     -- Stage 57
     -- Stage 58
     -- Stage 59
     -- Stage 60
     -- Stage 61
     -- Stage 62
     -- Stage 63
     -- Stage 64
     -- Stage 65
     -- Stage 66
     -- Stage 67
     -- Stage 68
     -- Stage 69
     -- Stage 70
     -- Stage 71
     -- Stage 72
     -- Stage 73
     -- Stage 74
     -- Stage 75
     -- Stage 76
     -- Stage 77
     -- Stage 78
     -- Stage 79
     -- Stage 80
     -- Stage 81
     -- Stage 82
     -- Stage 83
     -- Stage 84
     -- Stage 85
     -- Stage 86
     -- Stage 87
     -- Stage 88
     -- Stage 89
     -- Stage 90
     -- Stage 91
     -- Stage 92
     -- Stage 93
     -- Stage 94
     -- Stage 95
     -- Stage 96
     -- Stage 97
     -- Stage 98
     -- Stage 99
     -- Stage 100
     -- Stage 101
     -- Stage 102
     -- Stage 103
     -- Stage 104
     -- Stage 105
     -- Stage 106
     -- Stage 107
     -- Stage 108
     -- Stage 109
     -- Stage 110
     -- Stage 111
     -- Stage 112
     -- Stage 113
     -- Stage 114
     -- Stage 115
     -- Stage 116
     -- Stage 117
     -- Stage 118
     -- Stage 119
     -- Stage 120
     -- Stage 121
     -- Stage 122
     -- Stage 123
     -- Stage 124
     -- Stage 125
     -- Stage 126
     -- Stage 127
     -- Stage 128
     -- Stage 129
     -- Stage 130
     -- Stage 131
     -- Stage 132
     -- Stage 133
     -- Stage 134
     -- Stage 135
     -- Stage 136
     -- Stage 137
     -- Stage 138
     -- Stage 139
     -- Stage 140
     -- Stage 141
     -- Stage 142
     -- Stage 143
     -- Stage 144
     -- Stage 145
     -- Stage 146
     -- Stage 147
     -- Stage 148
     -- Stage 149
     -- Stage 150
     -- Stage 151
     -- Stage 152
     -- Stage 153
     -- Stage 154
     -- Stage 155
     -- Stage 156
     -- Stage 157
     -- Stage 158
     -- Stage 159
     -- Stage 160
     -- Stage 161
     -- Stage 162
     -- Stage 163
     -- Stage 164
     -- Stage 165
     -- Stage 166
     -- Stage 167
     -- Stage 168
     -- Stage 169
     -- Stage 170
     -- Stage 171
     -- Stage 172
     -- Stage 173
     -- Stage 174
     -- Stage 175
     -- Stage 176
     -- Stage 177
     -- Stage 178
     -- Stage 179
     -- Stage 180
     -- Stage 181
     -- Stage 182
     -- Stage 183
     -- Stage 184
     -- Stage 185
     -- Stage 186
     -- Stage 187
     -- Stage 188
     -- Stage 189
     -- Stage 190
     -- Stage 191
     -- Stage 192
     -- Stage 193
     -- Stage 194
     -- Stage 195
     -- Stage 196
     -- Stage 197
     -- Stage 198
     -- Stage 199
     -- Stage 200
     -- Stage 201
     -- Stage 202
     -- Stage 203
     -- Stage 204
     -- Stage 205
     -- Stage 206
     -- Stage 207
     -- Stage 208
     -- Stage 209
     -- Stage 210
     -- Stage 211
     -- Stage 212
     -- Stage 213
     -- Stage 214
     -- Stage 215
     -- Stage 216
     -- Stage 217
     -- Stage 218
     -- Stage 219
     -- Stage 220
     -- Stage 221
     -- Stage 222
     -- Stage 223
     -- Stage 224
     -- Stage 225
     -- Stage 226
     -- Stage 227
     -- Stage 228
     -- Stage 229
     -- Stage 230
     -- Stage 231
     -- Stage 232
     -- Stage 233
     -- Stage 234
     -- Stage 235
     -- Stage 236
     -- Stage 237
     -- Stage 238
     -- Stage 239
     -- Stage 240
     -- Stage 241
     -- Stage 242
     -- Stage 243
     -- Stage 244
     -- Stage 245
     -- Stage 246
     -- Stage 247
     -- Stage 248
     -- Stage 249
     -- Stage 250
     -- Stage 251
     -- Stage 252
     -- Stage 253
     -- Stage 254
     -- Stage 255
     -- Stage 256
     -- Stage 257
     -- Stage 258
     -- Stage 259
     -- Stage 260
     -- Stage 261
     -- Stage 262
     -- Stage 263
     -- Stage 264
     -- Stage 265
     -- Stage 266
     -- Stage 267
     -- Stage 268
     -- Stage 269
     -- Stage 270
     -- Stage 271
     -- Stage 272
     -- Stage 273
     -- Stage 274
     -- Stage 275
     -- Stage 276
     -- Stage 277
     -- Stage 278
     -- Stage 279
     -- Stage 280
     -- Stage 281
     -- Stage 282
     -- Stage 283
     -- Stage 284
     -- Stage 285
     -- Stage 286
     -- Stage 287
     -- Stage 288
     -- Stage 289
     -- Stage 290
     -- Stage 291
     -- Stage 292
     -- Stage 293
     -- Stage 294
     -- Stage 295
     -- Stage 296
     -- Stage 297
     -- Stage 298
     -- Stage 299
     -- Stage 300
     -- Stage 301
     -- Stage 302
     -- Stage 303
     -- Stage 304
     -- Stage 305
     -- Stage 306
     -- Stage 307
     -- Stage 308
     -- Stage 309
     -- Stage 310
     -- Stage 311
     -- Stage 312
     -- Stage 313
     -- Stage 314
     -- Stage 315
     -- Stage 316
     -- Stage 317
     -- Stage 318
     -- Stage 319
     -- Stage 320
     -- Stage 321
     -- Stage 322
     -- Stage 323
     -- Stage 324
     -- Stage 325
     -- Stage 326
     -- Stage 327
     -- Stage 328
     -- Stage 329
     -- Stage 330
     -- Stage 331
     -- Stage 332
     -- Stage 333
     -- Stage 334
     -- Stage 335
     -- Stage 336
     -- Stage 337
     -- Stage 338
     -- Stage 339
     -- Stage 340
     -- Stage 341
     -- Stage 342
     -- Stage 343
     -- Stage 344
     -- Stage 345
     -- Stage 346
     -- Stage 347
     -- Stage 348
     -- Stage 349
     -- Stage 350
     -- Stage 351
     -- Stage 352
     -- Stage 353
     -- Stage 354
     -- Stage 355
     -- Stage 356
     -- Stage 357
     -- Stage 358
     -- Stage 359
 end if;
end process;

end arch;
