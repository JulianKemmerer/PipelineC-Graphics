-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.001595949285482084, 0.012428088894585224, 0.023260228503688512, 0.03409236811279135, 0.044924507721894644, 0.05575664733099778, 0.06658878694010092, 0.07742092654920421, 0.08825306615830719, 0.09908520576741049, 0.10991734537651378, 0.12074948498561647, 0.1315816245947199, 0.14241376420382304, 0.1532459038129265, 0.16407804342202978, 0.17491018303113245, 0.18574232264023544, 0.19657446224933875, 0.20740660185844204, 0.21823874146754546, 0.22907088107664844, 0.23990302068575145, 0.2507351602948546, 0.261567299903958, 0.27239943951306084, 0.283231579122164, 0.29406371873126746, 0.3048958583403706, 0.3157279979494731, 0.32656013755857627, 0.3373922771676797, 0.3482244167767831, 0.35905655638588657, 0.3698886959949894, 0.38072083560409287, 0.3915529752131957, 0.40238511482229883, 0.41321725443140195, 0.4240493940405054, 0.43488153364960824, 0.445713673258712, 0.4565458128678148, 0.467377952476918, 0.4782100920860205, 0.48904223169512395, 0.49987437130422707, 0.5107065109133309, 0.5215386505224336, 0.5323707901315368, 0.5432029297406402, 0.5540350693497431, 0.5648672089588466, 0.5756993485679494, 0.5865314881770523, 0.5973636277861554, 0.6081957673952588, 0.6190279070043616, 0.6298600466134654, 0.6406921862225682, 0.6515243258316711, 0.6623564654407748, 0.6731886050498779, 0.6840207446589813, 0.6948528842680844, 0.705685023877187, 0.7165171634862905, 0.7273493030953939, 0.7381814427044965, 0.7490135823135996, 0.759845721922703, 0.7706778615318062, 0.781510001140909, 0.7923421407500124, 0.8031742803591162, 0.814006419968219, 0.8248385595773221, 0.8356706991864253, 0.8465028387955287, 0.8573349784046316, 0.8681671180137347, 0.8789992576228378, 0.8898313972319409, 0.9006635368410438, 0.911495676450147, 0.9223278160592504, 0.9331599556683535, 0.943992095277457, 0.9548242348865601, 0.9656563744956635, 0.9764885141047664, 0.9873206537138696, 0.9981527933229727]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 16
entity shade_183CLK_f33a2411 is
port(
 clk : in std_logic;
 global_to_module : in shade_global_to_module_t;
 background : in fixed3;
 dir : in float3;
 hit : in hit_out;
 hit_material : in material_t;
 minfog : in fixed;
 return_output : out fixed3);
end shade_183CLK_f33a2411;
architecture arch of shade_183CLK_f33a2411 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 183;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal REG_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal COMB_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 1
signal REG_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal REG_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal COMB_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 2
signal REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal REG_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal COMB_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 3
signal REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 4
signal REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 5
signal REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 6
signal REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 7
signal REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 8
signal REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 9
signal REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 10
signal REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 11
signal REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 12
signal REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 13
signal REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 14
signal REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 15
signal REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 16
signal REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 17
signal REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 18
signal REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 19
signal REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 20
signal REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 21
signal REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 22
signal REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 23
signal REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 24
signal REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 25
signal REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal REG_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
signal COMB_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
-- Stage 26
signal REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 27
signal REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 28
signal REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 29
signal REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 30
signal REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 31
signal REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 32
signal REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 33
signal REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 34
signal REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal REG_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal COMB_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 35
signal REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 36
signal REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 37
signal REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 38
signal REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 39
signal REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 40
signal REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 41
signal REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 42
signal REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 43
signal REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 44
signal REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 45
signal REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 46
signal REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 47
signal REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 48
signal REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 49
signal REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 50
signal REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 51
signal REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 52
signal REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 53
signal REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 54
signal REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 55
signal REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 56
signal REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 57
signal REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 58
signal REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 59
signal REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 60
signal REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 61
signal REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 62
signal REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 63
signal REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 64
signal REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 65
signal REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 66
signal REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 67
signal REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 68
signal REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 69
signal REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 70
signal REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 71
signal REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 72
signal REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 73
signal REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 74
signal REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 75
signal REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 76
signal REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 77
signal REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 78
signal REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 79
signal REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 80
signal REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 81
signal REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 82
signal REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 83
signal REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 84
signal REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 85
signal REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 86
signal REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 87
signal REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 88
signal REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 89
signal REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 90
signal REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 91
signal REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 92
signal REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 93
signal REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 94
signal REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 95
signal REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 96
signal REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 97
signal REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 98
signal REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 99
signal REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 100
signal REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 101
signal REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 102
signal REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 103
signal REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 104
signal REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 105
signal REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 106
signal REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 107
signal REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 108
signal REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 109
signal REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 110
signal REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 111
signal REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 112
signal REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 113
signal REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 114
signal REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 115
signal REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 116
signal REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 117
signal REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 118
signal REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 119
signal REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 120
signal REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 121
signal REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 122
signal REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 123
signal REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 124
signal REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 125
signal REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 126
signal REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 127
signal REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 128
signal REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 129
signal REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 130
signal REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 131
signal REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 132
signal REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 133
signal REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 134
signal REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 135
signal REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 136
signal REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 137
signal REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 138
signal REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 139
signal REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 140
signal REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 141
signal REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 142
signal REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 143
signal REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 144
signal REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 145
signal REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 146
signal REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 147
signal REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 148
signal REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 149
signal REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 150
signal REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 151
signal REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 152
signal REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 153
signal REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 154
signal REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 155
signal REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 156
signal REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 157
signal REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 158
signal REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 159
signal REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 160
signal REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 161
signal REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 162
signal REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 163
signal REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 164
signal REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 165
signal REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 166
signal REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 167
signal REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 168
signal REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 169
signal REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 170
signal REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal REG_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal COMB_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 171
signal REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 172
signal REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 173
signal REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 174
signal REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 175
signal REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal REG_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal REG_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal COMB_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal COMB_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
-- Stage 176
signal REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
-- Stage 177
signal REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
-- Stage 178
signal REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
-- Stage 179
signal REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
-- Stage 180
signal REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
-- Stage 181
signal REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal COMB_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal COMB_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
-- Stage 182
-- Each function instance gets signals
-- scene_colors[tr_pipelinec_gen_c_l370_c27_588d]
signal scene_colors_tr_pipelinec_gen_c_l370_c27_588d_scene : scene_t;
signal scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output : scene_colors_t;

-- BIN_OP_SL[tr_pipelinec_gen_c_l372_c27_7020]
signal BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_left : std_logic_vector(22 downto 0);
signal BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_right : signed(4 downto 0);
signal BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output : std_logic_vector(22 downto 0);

-- BIN_OP_LT[tr_pipelinec_gen_c_l374_c6_5562]
signal BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_left : std_logic_vector(22 downto 0);
signal BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_right : std_logic_vector(22 downto 0);
signal BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output : unsigned(0 downto 0);

-- rcolor_MUX[tr_pipelinec_gen_c_l374_c3_c373]
signal rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
signal rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iftrue : fixed3;
signal rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
signal rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output : fixed3;

-- reflect[tr_pipelinec_gen_c_l377_c22_9032]
signal reflect_tr_pipelinec_gen_c_l377_c22_9032_I : float3;
signal reflect_tr_pipelinec_gen_c_l377_c22_9032_N : float3;
signal reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output : float3;

-- cast_ray_nested[tr_pipelinec_gen_c_l378_c28_f218]
signal cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_hitin : point_and_dir;
signal cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output : fixed3;

-- light_intensity[tr_pipelinec_gen_c_l379_c16_e83f]
signal light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_hit : float3;
signal light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output : fixed;

-- fixed_make_from_double[tr_pipelinec_gen_c_l380_c88_ab10]
signal fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_a : std_logic_vector(22 downto 0);
signal fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output : fixed;

-- fixed_add[tr_pipelinec_gen_c_l380_c74_e9ac]
signal fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_left : fixed;
signal fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_right : fixed;
signal fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output : fixed;

-- fixed3_mul_fixed[tr_pipelinec_gen_c_l380_c28_2752]
signal fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
signal fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_right : fixed;
signal fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output : fixed3;

-- fixed3_mul[tr_pipelinec_gen_c_l381_c51_a739]
signal fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_left : fixed3;
signal fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
signal fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output : fixed3;

-- fixed3_add[tr_pipelinec_gen_c_l381_c25_97f1]
signal fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
signal fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_right : fixed3;
signal fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output : fixed3;

-- fixed_make_from_float[tr_pipelinec_gen_c_l382_c37_b99d]
signal fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_a : std_logic_vector(22 downto 0);
signal fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output : fixed;

-- color_max[tr_pipelinec_gen_c_l382_c27_3728]
signal color_max_tr_pipelinec_gen_c_l382_c27_3728_a : fixed;
signal color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
signal color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output : fixed;

-- color_select[tr_pipelinec_gen_c_l382_c14_e64f]
signal color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
signal color_select_tr_pipelinec_gen_c_l382_c14_e64f_a : fixed3;
signal color_select_tr_pipelinec_gen_c_l382_c14_e64f_b : fixed3;
signal color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output : fixed3;

function CONST_REF_RD_point_and_dir_point_and_dir_8057( ref_toks_0 : float3;
 ref_toks_1 : float3) return point_and_dir is
 
  variable base : point_and_dir; 
  variable return_output : point_and_dir;
begin
      base.orig := ref_toks_0;
      base.dir := ref_toks_1;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- scene_colors_tr_pipelinec_gen_c_l370_c27_588d
scene_colors_tr_pipelinec_gen_c_l370_c27_588d : entity work.scene_colors_0CLK_5af1a430 port map (
scene_colors_tr_pipelinec_gen_c_l370_c27_588d_scene,
scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output);

-- BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020
BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020 : entity work.BIN_OP_SL_float_8_14_t_int5_t_1CLK_9d8547c8 port map (
clk,
BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_left,
BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_right,
BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output);

-- BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562
BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562 : entity work.BIN_OP_LT_float_8_14_t_float_8_14_t_1CLK_6a161d44 port map (
clk,
BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_left,
BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_right,
BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output);

-- rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373
rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373 : entity work.MUX_uint1_t_fixed3_fixed3_1CLK_dafad20f port map (
clk,
rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iftrue,
rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output);

-- reflect_tr_pipelinec_gen_c_l377_c22_9032
reflect_tr_pipelinec_gen_c_l377_c22_9032 : entity work.reflect_26CLK_48b4560d port map (
clk,
reflect_tr_pipelinec_gen_c_l377_c22_9032_I,
reflect_tr_pipelinec_gen_c_l377_c22_9032_N,
reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output);

-- cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218
cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218 : entity work.cast_ray_nested_145CLK_96264b07 port map (
clk,
global_to_module.cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218,
cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_hitin,
cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output);

-- light_intensity_tr_pipelinec_gen_c_l379_c16_e83f
light_intensity_tr_pipelinec_gen_c_l379_c16_e83f : entity work.light_intensity_34CLK_55880f91 port map (
clk,
light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_hit,
light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output);

-- fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10
fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10 : entity work.fixed_make_from_double_0CLK_38477f9e port map (
fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_a,
fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output);

-- fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac
fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac : entity work.fixed_add_1CLK_419e1dd2 port map (
clk,
fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_left,
fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_right,
fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output);

-- fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752
fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752 : entity work.fixed3_mul_fixed_5CLK_c4855664 port map (
clk,
fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_right,
fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output);

-- fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739
fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739 : entity work.fixed3_mul_5CLK_40e12b03 port map (
clk,
fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_left,
fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output);

-- fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1
fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1 : entity work.fixed3_add_0CLK_f982eca9 port map (
fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_right,
fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output);

-- fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d
fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d : entity work.fixed_make_from_float_2CLK_c0caf0ba port map (
clk,
fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_a,
fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output);

-- color_max_tr_pipelinec_gen_c_l382_c27_3728
color_max_tr_pipelinec_gen_c_l382_c27_3728 : entity work.color_max_1CLK_71e85ea2 port map (
clk,
color_max_tr_pipelinec_gen_c_l382_c27_3728_a,
color_max_tr_pipelinec_gen_c_l382_c27_3728_b,
color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output);

-- color_select_tr_pipelinec_gen_c_l382_c14_e64f
color_select_tr_pipelinec_gen_c_l382_c14_e64f : entity work.color_select_6CLK_94dcec9d port map (
clk,
color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
color_select_tr_pipelinec_gen_c_l382_c14_e64f_a,
color_select_tr_pipelinec_gen_c_l382_c14_e64f_b,
color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 background,
 dir,
 hit,
 hit_material,
 minfog,
 -- Registers
 -- Stage 0
 REG_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b,
 REG_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 1
 REG_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b,
 REG_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 2
 REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b,
 REG_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 3
 REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 4
 REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 5
 REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 6
 REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 7
 REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 8
 REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 9
 REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 10
 REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 11
 REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 12
 REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 13
 REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 14
 REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 15
 REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 16
 REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 17
 REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 18
 REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 19
 REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 20
 REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 21
 REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 22
 REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 23
 REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 24
 REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 25
 REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 REG_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
 -- Stage 26
 REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 27
 REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 28
 REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 29
 REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 30
 REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 31
 REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 32
 REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 33
 REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 34
 REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left,
 REG_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 35
 REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 36
 REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 37
 REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 38
 REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 39
 REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 40
 REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 41
 REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 42
 REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 43
 REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 44
 REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 45
 REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 46
 REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 47
 REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 48
 REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 49
 REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 50
 REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 51
 REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 52
 REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 53
 REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 54
 REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 55
 REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 56
 REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 57
 REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 58
 REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 59
 REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 60
 REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 61
 REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 62
 REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 63
 REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 64
 REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 65
 REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 66
 REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 67
 REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 68
 REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 69
 REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 70
 REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 71
 REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 72
 REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 73
 REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 74
 REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 75
 REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 76
 REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 77
 REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 78
 REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 79
 REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 80
 REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 81
 REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 82
 REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 83
 REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 84
 REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 85
 REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 86
 REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 87
 REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 88
 REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 89
 REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 90
 REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 91
 REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 92
 REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 93
 REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 94
 REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 95
 REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 96
 REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 97
 REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 98
 REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 99
 REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 100
 REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 101
 REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 102
 REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 103
 REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 104
 REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 105
 REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 106
 REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 107
 REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 108
 REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 109
 REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 110
 REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 111
 REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 112
 REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 113
 REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 114
 REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 115
 REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 116
 REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 117
 REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 118
 REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 119
 REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 120
 REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 121
 REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 122
 REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 123
 REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 124
 REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 125
 REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 126
 REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 127
 REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 128
 REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 129
 REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 130
 REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 131
 REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 132
 REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 133
 REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 134
 REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 135
 REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 136
 REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 137
 REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 138
 REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 139
 REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 140
 REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 141
 REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 142
 REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 143
 REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 144
 REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 145
 REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 146
 REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 147
 REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 148
 REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 149
 REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 150
 REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 151
 REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 152
 REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 153
 REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 154
 REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 155
 REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 156
 REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 157
 REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 158
 REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 159
 REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 160
 REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 161
 REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 162
 REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 163
 REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 164
 REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 165
 REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 166
 REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 167
 REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 168
 REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 169
 REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 170
 REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right,
 REG_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 171
 REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 172
 REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 173
 REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 174
 REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 175
 REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 REG_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left,
 REG_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x,
 -- Stage 176
 REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 -- Stage 177
 REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 -- Stage 178
 REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 -- Stage 179
 REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 -- Stage 180
 REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 -- Stage 181
 REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse,
 REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond,
 -- Stage 182
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output,
 BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output,
 BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output,
 rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output,
 reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output,
 cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output,
 light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output,
 fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output,
 fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output,
 fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output,
 fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output,
 fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output,
 fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output,
 color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output,
 color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : fixed3;
 variable VAR_background : fixed3;
 variable VAR_dir : float3;
 variable VAR_hit : hit_out;
 variable VAR_hit_material : material_t;
 variable VAR_minfog : fixed;
 variable VAR_state : full_state_t;
 variable VAR_scene : scene_t;
 variable VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l369_c19_7d7e_return_output : scene_t;
 variable VAR_colors : scene_colors_t;
 variable VAR_scene_colors_tr_pipelinec_gen_c_l370_c27_588d_scene : scene_t;
 variable VAR_scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output : scene_colors_t;
 variable VAR_rcolor : fixed3;
 variable VAR_fogmix : std_logic_vector(22 downto 0);
 variable VAR_CONST_REF_RD_float_8_14_t_hit_out_dist_d41d_tr_pipelinec_gen_c_l372_c27_bc68_return_output : std_logic_vector(22 downto 0);
 variable VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_left : std_logic_vector(22 downto 0);
 variable VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_right : signed(4 downto 0);
 variable VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output : std_logic_vector(22 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_left : std_logic_vector(22 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_right : std_logic_vector(22 downto 0);
 variable VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output : unsigned(0 downto 0);
 variable VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iftrue : fixed3;
 variable VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse : fixed3;
 variable VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output : fixed3;
 variable VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond : unsigned(0 downto 0);
 variable VAR_hitreflect : point_and_dir;
 variable VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_I : float3;
 variable VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_N : float3;
 variable VAR_CONST_REF_RD_float3_hit_out_hit_dir_d41d_tr_pipelinec_gen_c_l377_c35_3513_return_output : float3;
 variable VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output : float3;
 variable VAR_reflect_color : fixed3;
 variable VAR_cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_hitin : point_and_dir;
 variable VAR_CONST_REF_RD_point_and_dir_point_and_dir_8057_tr_pipelinec_gen_c_l378_c44_0f5e_return_output : point_and_dir;
 variable VAR_cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output : fixed3;
 variable VAR_li : fixed;
 variable VAR_light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_hit : float3;
 variable VAR_light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output : fixed;
 variable VAR_diffuse_color : fixed3;
 variable VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left : fixed3;
 variable VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_right : fixed;
 variable VAR_CONST_REF_RD_fixed3_material_t_diffuse_color_d41d_tr_pipelinec_gen_c_l380_c45_eded_return_output : fixed3;
 variable VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_left : fixed;
 variable VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_right : fixed;
 variable VAR_fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_a : std_logic_vector(22 downto 0);
 variable VAR_fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output : fixed;
 variable VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output : fixed;
 variable VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output : fixed3;
 variable VAR_comb_color : fixed3;
 variable VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left : fixed3;
 variable VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_right : fixed3;
 variable VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_left : fixed3;
 variable VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right : fixed3;
 variable VAR_CONST_REF_RD_fixed3_material_t_reflect_color_d41d_tr_pipelinec_gen_c_l381_c77_abf0_return_output : fixed3;
 variable VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output : fixed3;
 variable VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output : fixed3;
 variable VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x : fixed;
 variable VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_a : fixed3;
 variable VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_b : fixed3;
 variable VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_a : fixed;
 variable VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b : fixed;
 variable VAR_fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_a : std_logic_vector(22 downto 0);
 variable VAR_fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output : fixed;
 variable VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output : fixed;
 variable VAR_CONST_REF_RD_fixed3_scene_colors_t_fog_d41d_tr_pipelinec_gen_c_l382_c77_b397_return_output : fixed3;
 variable VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output : fixed3;
 variable VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output : float3;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_a := to_slv(to_float(0.2, 8, 14));
     VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_right := to_signed(-9, 5);
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_right := to_slv(to_float(1.0, 8, 14));
     -- fixed_make_from_double[tr_pipelinec_gen_c_l380_c88_ab10] LATENCY=0
     -- Inputs
     fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_a <= VAR_fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_a;
     -- Outputs
     VAR_fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output := fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output;

     -- Submodule level 1
     VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_right := VAR_fixed_make_from_double_tr_pipelinec_gen_c_l380_c88_ab10_return_output;
 -- Reads from global variables
     VAR_state := global_to_module.state;
     -- Submodule level 0
     -- CONST_REF_RD_scene_t_full_state_t_scene_d41d[tr_pipelinec_gen_c_l369_c19_7d7e] LATENCY=0
     VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l369_c19_7d7e_return_output := VAR_state.scene;

     -- Submodule level 1
     VAR_scene_colors_tr_pipelinec_gen_c_l370_c27_588d_scene := VAR_CONST_REF_RD_scene_t_full_state_t_scene_d41d_tr_pipelinec_gen_c_l369_c19_7d7e_return_output;
     -- scene_colors[tr_pipelinec_gen_c_l370_c27_588d] LATENCY=0
     -- Inputs
     scene_colors_tr_pipelinec_gen_c_l370_c27_588d_scene <= VAR_scene_colors_tr_pipelinec_gen_c_l370_c27_588d_scene;
     -- Outputs
     VAR_scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output := scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_fixed3_scene_colors_t_fog_d41d[tr_pipelinec_gen_c_l382_c77_b397] LATENCY=0
     VAR_CONST_REF_RD_fixed3_scene_colors_t_fog_d41d_tr_pipelinec_gen_c_l382_c77_b397_return_output := VAR_scene_colors_tr_pipelinec_gen_c_l370_c27_588d_return_output.fog;

     -- Submodule level 3
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_a := VAR_CONST_REF_RD_fixed3_scene_colors_t_fog_d41d_tr_pipelinec_gen_c_l382_c77_b397_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_background := background;
     VAR_dir := dir;
     VAR_hit := hit;
     VAR_hit_material := hit_material;
     VAR_minfog := minfog;

     -- Submodule level 0
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := VAR_background;
     VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_I := VAR_dir;
     VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b := VAR_minfog;
     -- CONST_REF_RD_float_8_14_t_hit_out_dist_d41d[tr_pipelinec_gen_c_l372_c27_bc68] LATENCY=0
     VAR_CONST_REF_RD_float_8_14_t_hit_out_dist_d41d_tr_pipelinec_gen_c_l372_c27_bc68_return_output := VAR_hit.dist;

     -- CONST_REF_RD_float3_hit_out_hit_dir_d41d[tr_pipelinec_gen_c_l377_c35_3513] LATENCY=0
     VAR_CONST_REF_RD_float3_hit_out_hit_dir_d41d_tr_pipelinec_gen_c_l377_c35_3513_return_output := VAR_hit.hit.dir;

     -- CONST_REF_RD_fixed3_material_t_reflect_color_d41d[tr_pipelinec_gen_c_l381_c77_abf0] LATENCY=0
     VAR_CONST_REF_RD_fixed3_material_t_reflect_color_d41d_tr_pipelinec_gen_c_l381_c77_abf0_return_output := VAR_hit_material.reflect_color;

     -- CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f LATENCY=0
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := VAR_hit.hit.orig;

     -- CONST_REF_RD_fixed3_material_t_diffuse_color_d41d[tr_pipelinec_gen_c_l380_c45_eded] LATENCY=0
     VAR_CONST_REF_RD_fixed3_material_t_diffuse_color_d41d_tr_pipelinec_gen_c_l380_c45_eded_return_output := VAR_hit_material.diffuse_color;

     -- Submodule level 1
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := VAR_CONST_REF_RD_fixed3_material_t_diffuse_color_d41d_tr_pipelinec_gen_c_l380_c45_eded_return_output;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := VAR_CONST_REF_RD_fixed3_material_t_reflect_color_d41d_tr_pipelinec_gen_c_l381_c77_abf0_return_output;
     VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_N := VAR_CONST_REF_RD_float3_hit_out_hit_dir_d41d_tr_pipelinec_gen_c_l377_c35_3513_return_output;
     VAR_light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_hit := VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_left := VAR_CONST_REF_RD_float_8_14_t_hit_out_dist_d41d_tr_pipelinec_gen_c_l372_c27_bc68_return_output;
     -- BIN_OP_SL[tr_pipelinec_gen_c_l372_c27_7020] LATENCY=1
     -- Inputs
     BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_left <= VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_left;
     BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_right <= VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_right;

     -- light_intensity[tr_pipelinec_gen_c_l379_c16_e83f] LATENCY=34
     -- Inputs
     light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_hit <= VAR_light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_hit;

     -- reflect[tr_pipelinec_gen_c_l377_c22_9032] LATENCY=26
     -- Inputs
     reflect_tr_pipelinec_gen_c_l377_c22_9032_I <= VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_I;
     reflect_tr_pipelinec_gen_c_l377_c22_9032_N <= VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_N;

     -- Write to comb signals
     COMB_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     COMB_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b := REG_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Submodule outputs
     VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output := BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output;

     -- Submodule level 0
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_left := VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output;
     VAR_fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_a := VAR_BIN_OP_SL_tr_pipelinec_gen_c_l372_c27_7020_return_output;
     -- BIN_OP_LT[tr_pipelinec_gen_c_l374_c6_5562] LATENCY=1
     -- Inputs
     BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_left <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_left;
     BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_right <= VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_right;

     -- fixed_make_from_float[tr_pipelinec_gen_c_l382_c37_b99d] LATENCY=2
     -- Inputs
     fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_a <= VAR_fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_a;

     -- Write to comb signals
     COMB_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     COMB_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b := REG_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Submodule outputs
     VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output := BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output;

     -- Submodule level 0
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := VAR_BIN_OP_LT_tr_pipelinec_gen_c_l374_c6_5562_return_output;
     -- Write to comb signals
     COMB_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     COMB_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b := REG_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Submodule outputs
     VAR_fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output := fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output;

     -- Submodule level 0
     VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_a := VAR_fixed_make_from_float_tr_pipelinec_gen_c_l382_c37_b99d_return_output;
     -- color_max[tr_pipelinec_gen_c_l382_c27_3728] LATENCY=1
     -- Inputs
     color_max_tr_pipelinec_gen_c_l382_c27_3728_a <= VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_a;
     color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;

     -- Write to comb signals
     COMB_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Submodule outputs
     VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output := color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output;

     -- Submodule level 0
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := VAR_color_max_tr_pipelinec_gen_c_l382_c27_3728_return_output;
     -- Write to comb signals
     COMB_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 7 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 13 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 14 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 15 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 16 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 17 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 18 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 19 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 20 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 21 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 22 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 23 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 24 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 25 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;

     -- Write to comb signals
     COMB_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     COMB_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
   elsif STAGE = 26 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output := REG_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Submodule outputs
     VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output := reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output;

     -- Submodule level 0
     -- CONST_REF_RD_point_and_dir_point_and_dir_8057[tr_pipelinec_gen_c_l378_c44_0f5e] LATENCY=0
     VAR_CONST_REF_RD_point_and_dir_point_and_dir_8057_tr_pipelinec_gen_c_l378_c44_0f5e_return_output := CONST_REF_RD_point_and_dir_point_and_dir_8057(
     VAR_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output,
     VAR_reflect_tr_pipelinec_gen_c_l377_c22_9032_return_output);

     -- Submodule level 1
     VAR_cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_hitin := VAR_CONST_REF_RD_point_and_dir_point_and_dir_8057_tr_pipelinec_gen_c_l378_c44_0f5e_return_output;
     -- cast_ray_nested[tr_pipelinec_gen_c_l378_c28_f218] LATENCY=145
     -- Inputs
     cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_hitin <= VAR_cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_hitin;

     -- Write to comb signals
     COMB_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 27 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 28 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 29 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 30 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 31 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 32 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 33 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 34 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Submodule outputs
     VAR_light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output := light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output;

     -- Submodule level 0
     VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_left := VAR_light_intensity_tr_pipelinec_gen_c_l379_c16_e83f_return_output;
     -- fixed_add[tr_pipelinec_gen_c_l380_c74_e9ac] LATENCY=1
     -- Inputs
     fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_left <= VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_left;
     fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_right <= VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_right;

     -- Write to comb signals
     COMB_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     COMB_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 35 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left := REG_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Submodule outputs
     VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output := fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output;

     -- Submodule level 0
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_right := VAR_fixed_add_tr_pipelinec_gen_c_l380_c74_e9ac_return_output;
     -- fixed3_mul_fixed[tr_pipelinec_gen_c_l380_c28_2752] LATENCY=5
     -- Inputs
     fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_right <= VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_right;

     -- Write to comb signals
     COMB_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 36 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 37 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 38 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 39 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 40 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Submodule outputs
     VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output := fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output;

     -- Submodule level 0
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := VAR_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_return_output;
     -- Write to comb signals
     COMB_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 41 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 42 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 43 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 44 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 45 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 46 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 47 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 48 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 49 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 50 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 51 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 52 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 53 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 54 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 55 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 56 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 57 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 58 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 59 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 60 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 61 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 62 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 63 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 64 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 65 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 66 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 67 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 68 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 69 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 70 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 71 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 72 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 73 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 74 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 75 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 76 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 77 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 78 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 79 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 80 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 81 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 82 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 83 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 84 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 85 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 86 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 87 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 88 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 89 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 90 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 91 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 92 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 93 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 94 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 95 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 96 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 97 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 98 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 99 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 100 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 101 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 102 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 103 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 104 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 105 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 106 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 107 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 108 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 109 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 110 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 111 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 112 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 113 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 114 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 115 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 116 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 117 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 118 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 119 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 120 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 121 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 122 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 123 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 124 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 125 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 126 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 127 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 128 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 129 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 130 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 131 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 132 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 133 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 134 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 135 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 136 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 137 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 138 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 139 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 140 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 141 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 142 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 143 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 144 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 145 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 146 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 147 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 148 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 149 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 150 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 151 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 152 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 153 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 154 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 155 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 156 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 157 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 158 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 159 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 160 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 161 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 162 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 163 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 164 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 165 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 166 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 167 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 168 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 169 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 170 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     COMB_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 171 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right := REG_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Submodule outputs
     VAR_cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output := cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output;

     -- Submodule level 0
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_left := VAR_cast_ray_nested_tr_pipelinec_gen_c_l378_c28_f218_return_output;
     -- fixed3_mul[tr_pipelinec_gen_c_l381_c51_a739] LATENCY=5
     -- Inputs
     fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_left <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_left;
     fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;

     -- Write to comb signals
     COMB_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 172 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 173 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 174 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 175 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;

     -- Write to comb signals
     COMB_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     COMB_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     COMB_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
   elsif STAGE = 176 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left := REG_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x := REG_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Submodule outputs
     VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output := fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output;

     -- Submodule level 0
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_right := VAR_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_return_output;
     -- fixed3_add[tr_pipelinec_gen_c_l381_c25_97f1] LATENCY=0
     -- Inputs
     fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_right <= VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_right;
     -- Outputs
     VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output := fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output;

     -- Submodule level 1
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_b := VAR_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_return_output;
     -- color_select[tr_pipelinec_gen_c_l382_c14_e64f] LATENCY=6
     -- Inputs
     color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     color_select_tr_pipelinec_gen_c_l382_c14_e64f_a <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_a;
     color_select_tr_pipelinec_gen_c_l382_c14_e64f_b <= VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_b;

     -- Write to comb signals
     COMB_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
   elsif STAGE = 177 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;

     -- Write to comb signals
     COMB_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
   elsif STAGE = 178 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;

     -- Write to comb signals
     COMB_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
   elsif STAGE = 179 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;

     -- Write to comb signals
     COMB_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
   elsif STAGE = 180 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;

     -- Write to comb signals
     COMB_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
   elsif STAGE = 181 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;

     -- Write to comb signals
     COMB_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     COMB_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
   elsif STAGE = 182 then
     -- Read from prev stage
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse := REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond := REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Submodule outputs
     VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output := color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output;

     -- Submodule level 0
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iftrue := VAR_color_select_tr_pipelinec_gen_c_l382_c14_e64f_return_output;
     -- rcolor_MUX[tr_pipelinec_gen_c_l374_c3_c373] LATENCY=1
     -- Inputs
     rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iftrue <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iftrue;
     rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;

     -- Write to comb signals
   elsif STAGE = 183 then
     -- Read from prev stage
     -- Submodule outputs
     VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output := rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output;

     -- Submodule level 0
     VAR_return_output := VAR_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
     -- Stage 0
     REG_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE0_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE0_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE0_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= COMB_STAGE0_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     REG_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE0_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 1
     REG_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE1_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE1_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE1_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= COMB_STAGE1_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     REG_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE1_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 2
     REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE2_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE2_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE2_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b <= COMB_STAGE2_color_max_tr_pipelinec_gen_c_l382_c27_3728_b;
     REG_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE2_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 3
     REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE3_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE3_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE3_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE3_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 4
     REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE4_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE4_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE4_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE4_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE4_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 5
     REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE5_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE5_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE5_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE5_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE5_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 6
     REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE6_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE6_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE6_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE6_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE6_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 7
     REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE7_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE7_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE7_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE7_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE7_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 8
     REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE8_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE8_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE8_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE8_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE8_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 9
     REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE9_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE9_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE9_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE9_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE9_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 10
     REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE10_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE10_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE10_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE10_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE10_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 11
     REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE11_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE11_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE11_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE11_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE11_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 12
     REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE12_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE12_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE12_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE12_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE12_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 13
     REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE13_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE13_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE13_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE13_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE13_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 14
     REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE14_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE14_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE14_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE14_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE14_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 15
     REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE15_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE15_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE15_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE15_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE15_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 16
     REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE16_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE16_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE16_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE16_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE16_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 17
     REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE17_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE17_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE17_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE17_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE17_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 18
     REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE18_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE18_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE18_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE18_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE18_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 19
     REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE19_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE19_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE19_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE19_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE19_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 20
     REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE20_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE20_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE20_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE20_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE20_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 21
     REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE21_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE21_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE21_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE21_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE21_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 22
     REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE22_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE22_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE22_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE22_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE22_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 23
     REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE23_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE23_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE23_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE23_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE23_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 24
     REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE24_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE24_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE24_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE24_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE24_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 25
     REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE25_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE25_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE25_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE25_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     REG_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output <= COMB_STAGE25_CONST_REF_RD_float3_hit_out_hit_orig_d41d_tr_pipelinec_gen_c_l379_l376_DUPLICATE_e82f_return_output;
     -- Stage 26
     REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE26_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE26_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE26_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE26_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 27
     REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE27_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE27_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE27_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE27_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 28
     REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE28_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE28_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE28_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE28_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 29
     REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE29_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE29_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE29_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE29_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 30
     REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE30_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE30_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE30_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE30_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 31
     REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE31_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE31_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE31_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE31_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 32
     REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE32_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE32_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE32_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE32_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 33
     REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE33_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE33_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE33_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE33_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 34
     REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE34_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left <= COMB_STAGE34_fixed3_mul_fixed_tr_pipelinec_gen_c_l380_c28_2752_left;
     REG_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE34_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE34_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 35
     REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE35_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE35_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE35_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 36
     REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE36_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE36_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE36_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 37
     REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE37_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE37_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE37_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 38
     REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE38_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE38_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE38_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 39
     REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE39_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE39_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE39_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 40
     REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE40_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE40_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE40_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE40_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 41
     REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE41_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE41_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE41_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE41_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 42
     REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE42_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE42_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE42_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE42_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 43
     REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE43_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE43_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE43_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE43_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 44
     REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE44_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE44_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE44_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE44_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 45
     REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE45_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE45_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE45_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE45_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 46
     REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE46_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE46_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE46_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE46_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 47
     REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE47_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE47_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE47_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE47_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 48
     REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE48_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE48_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE48_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE48_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 49
     REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE49_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE49_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE49_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE49_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 50
     REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE50_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE50_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE50_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE50_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 51
     REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE51_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE51_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE51_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE51_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 52
     REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE52_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE52_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE52_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE52_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 53
     REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE53_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE53_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE53_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE53_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 54
     REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE54_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE54_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE54_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE54_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 55
     REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE55_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE55_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE55_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE55_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 56
     REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE56_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE56_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE56_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE56_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 57
     REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE57_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE57_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE57_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE57_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 58
     REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE58_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE58_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE58_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE58_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 59
     REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE59_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE59_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE59_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE59_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 60
     REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE60_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE60_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE60_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE60_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 61
     REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE61_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE61_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE61_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE61_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 62
     REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE62_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE62_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE62_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE62_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 63
     REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE63_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE63_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE63_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE63_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 64
     REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE64_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE64_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE64_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE64_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 65
     REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE65_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE65_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE65_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE65_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 66
     REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE66_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE66_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE66_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE66_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 67
     REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE67_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE67_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE67_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE67_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 68
     REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE68_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE68_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE68_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE68_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 69
     REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE69_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE69_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE69_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE69_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 70
     REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE70_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE70_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE70_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE70_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 71
     REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE71_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE71_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE71_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE71_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 72
     REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE72_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE72_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE72_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE72_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 73
     REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE73_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE73_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE73_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE73_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 74
     REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE74_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE74_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE74_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE74_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 75
     REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE75_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE75_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE75_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE75_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 76
     REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE76_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE76_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE76_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE76_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 77
     REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE77_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE77_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE77_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE77_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 78
     REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE78_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE78_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE78_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE78_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 79
     REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE79_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE79_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE79_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE79_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 80
     REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE80_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE80_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE80_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE80_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 81
     REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE81_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE81_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE81_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE81_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 82
     REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE82_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE82_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE82_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE82_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 83
     REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE83_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE83_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE83_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE83_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 84
     REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE84_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE84_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE84_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE84_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 85
     REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE85_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE85_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE85_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE85_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 86
     REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE86_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE86_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE86_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE86_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 87
     REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE87_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE87_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE87_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE87_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 88
     REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE88_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE88_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE88_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE88_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 89
     REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE89_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE89_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE89_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE89_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 90
     REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE90_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE90_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE90_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE90_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 91
     REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE91_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE91_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE91_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE91_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 92
     REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE92_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE92_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE92_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE92_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 93
     REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE93_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE93_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE93_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE93_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 94
     REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE94_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE94_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE94_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE94_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 95
     REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE95_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE95_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE95_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE95_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 96
     REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE96_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE96_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE96_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE96_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 97
     REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE97_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE97_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE97_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE97_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 98
     REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE98_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE98_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE98_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE98_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 99
     REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE99_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE99_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE99_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE99_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 100
     REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE100_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE100_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE100_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE100_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 101
     REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE101_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE101_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE101_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE101_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 102
     REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE102_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE102_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE102_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE102_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 103
     REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE103_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE103_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE103_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE103_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 104
     REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE104_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE104_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE104_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE104_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 105
     REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE105_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE105_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE105_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE105_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 106
     REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE106_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE106_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE106_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE106_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 107
     REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE107_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE107_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE107_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE107_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 108
     REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE108_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE108_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE108_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE108_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 109
     REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE109_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE109_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE109_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE109_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 110
     REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE110_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE110_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE110_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE110_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 111
     REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE111_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE111_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE111_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE111_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 112
     REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE112_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE112_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE112_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE112_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 113
     REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE113_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE113_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE113_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE113_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 114
     REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE114_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE114_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE114_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE114_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 115
     REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE115_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE115_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE115_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE115_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 116
     REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE116_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE116_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE116_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE116_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 117
     REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE117_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE117_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE117_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE117_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 118
     REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE118_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE118_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE118_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE118_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 119
     REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE119_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE119_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE119_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE119_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 120
     REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE120_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE120_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE120_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE120_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 121
     REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE121_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE121_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE121_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE121_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 122
     REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE122_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE122_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE122_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE122_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 123
     REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE123_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE123_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE123_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE123_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 124
     REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE124_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE124_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE124_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE124_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 125
     REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE125_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE125_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE125_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE125_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 126
     REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE126_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE126_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE126_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE126_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 127
     REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE127_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE127_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE127_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE127_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 128
     REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE128_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE128_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE128_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE128_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 129
     REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE129_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE129_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE129_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE129_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 130
     REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE130_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE130_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE130_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE130_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 131
     REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE131_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE131_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE131_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE131_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 132
     REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE132_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE132_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE132_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE132_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 133
     REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE133_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE133_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE133_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE133_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 134
     REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE134_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE134_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE134_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE134_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 135
     REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE135_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE135_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE135_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE135_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 136
     REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE136_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE136_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE136_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE136_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 137
     REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE137_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE137_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE137_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE137_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 138
     REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE138_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE138_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE138_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE138_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 139
     REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE139_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE139_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE139_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE139_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 140
     REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE140_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE140_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE140_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE140_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 141
     REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE141_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE141_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE141_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE141_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 142
     REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE142_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE142_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE142_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE142_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 143
     REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE143_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE143_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE143_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE143_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 144
     REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE144_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE144_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE144_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE144_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 145
     REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE145_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE145_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE145_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE145_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 146
     REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE146_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE146_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE146_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE146_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 147
     REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE147_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE147_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE147_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE147_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 148
     REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE148_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE148_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE148_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE148_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 149
     REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE149_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE149_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE149_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE149_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 150
     REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE150_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE150_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE150_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE150_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 151
     REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE151_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE151_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE151_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE151_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 152
     REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE152_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE152_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE152_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE152_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 153
     REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE153_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE153_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE153_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE153_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 154
     REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE154_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE154_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE154_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE154_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 155
     REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE155_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE155_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE155_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE155_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 156
     REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE156_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE156_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE156_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE156_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 157
     REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE157_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE157_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE157_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE157_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 158
     REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE158_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE158_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE158_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE158_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 159
     REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE159_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE159_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE159_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE159_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 160
     REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE160_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE160_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE160_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE160_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 161
     REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE161_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE161_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE161_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE161_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 162
     REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE162_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE162_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE162_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE162_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 163
     REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE163_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE163_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE163_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE163_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 164
     REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE164_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE164_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE164_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE164_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 165
     REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE165_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE165_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE165_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE165_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 166
     REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE166_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE166_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE166_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE166_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 167
     REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE167_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE167_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE167_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE167_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 168
     REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE168_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE168_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE168_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE168_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 169
     REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE169_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE169_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE169_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE169_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 170
     REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE170_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE170_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right <= COMB_STAGE170_fixed3_mul_tr_pipelinec_gen_c_l381_c51_a739_right;
     REG_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE170_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 171
     REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE171_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE171_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE171_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 172
     REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE172_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE172_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE172_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 173
     REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE173_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE173_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE173_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 174
     REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE174_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE174_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE174_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 175
     REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE175_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     REG_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left <= COMB_STAGE175_fixed3_add_tr_pipelinec_gen_c_l381_c25_97f1_left;
     REG_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x <= COMB_STAGE175_color_select_tr_pipelinec_gen_c_l382_c14_e64f_x;
     -- Stage 176
     REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE176_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Stage 177
     REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE177_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Stage 178
     REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE178_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Stage 179
     REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE179_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Stage 180
     REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE180_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Stage 181
     REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse <= COMB_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_iffalse;
     REG_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond <= COMB_STAGE181_rcolor_MUX_tr_pipelinec_gen_c_l374_c3_c373_cond;
     -- Stage 182
 end if;
end process;

end arch;
